magic
tech sky130A
timestamp 1618573301
<< xpolycontact >>
rect -201 -11 20 47
rect 510 -10 731 48
<< xpolyres >>
rect 20 0 510 35
<< end >>
