* SPICE3 file created from BGR.ext - technology: sky130A

.option scale=5000u

.subckt BGR GND Vref En
X0 E GND GND sky130_fd_pr__pnp_05v0 area=1.29416e+09
X1 A C w_16722_12162# w_16722_12162# sky130_fd_pr__pfet_g5v0d10v5 ad=72 pd=0 as=-1 ps=-1 w=4000 l=1000
X2 E GND GND sky130_fd_pr__pnp_05v0 area=0
X3 C C w_16722_12162# w_16722_12162# sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=-0 ps=-0 w=4000 l=1000
X4 E GND GND sky130_fd_pr__pnp_05v0 area=0
X5 E GND GND sky130_fd_pr__pnp_05v0 area=0
X6 H C w_16722_12162# w_16722_12162# sky130_fd_pr__pfet_g5v0d10v5 ad=113 pd=0 as=-0 ps=-0 w=4000 l=1000
X7 I GND GND sky130_fd_pr__pnp_05v0 area=1.27541e+09
X8 F GND GND sky130_fd_pr__pnp_05v0 area=113
X9 E GND GND sky130_fd_pr__pnp_05v0 area=0
X10 E GND GND sky130_fd_pr__pnp_05v0 area=0
X11 E GND GND sky130_fd_pr__pnp_05v0 area=0
X12 E GND GND sky130_fd_pr__pnp_05v0 area=0
X13 F Vref GND sky130_fd_pr__res_xhigh_po w=70 l=8720
X14 E J GND sky130_fd_pr__res_xhigh_po w=70 l=980
X15 w_16722_12162# K GND sky130_fd_pr__res_xhigh_po w=70 l=6924
X16 C G GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
X17 B En li_16144_1712# GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.29244e+09 pd=22081 as=897 ps=0 w=4000 l=1000
X18 A A B GND sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
X19 D A C GND sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
X20 J En D GND sky130_fd_pr__nfet_g5v0d10v5 ad=337 pd=0 as=0 ps=0 w=4000 l=1000
X21 Vref En H GND sky130_fd_pr__nfet_g5v0d10v5 ad=135 pd=0 as=0 ps=0 w=4000 l=1000
X22 K En G GND sky130_fd_pr__nfet_g5v0d10v5 ad=8 pd=0 as=8 ps=0 w=4000 l=1000
X23 G A GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=200
C0 li_16144_1712# J 1.02fF
C1 G C 0.06fF
C2 li_16144_1712# G 0.38fF
C3 Vref C 0.91fF
C4 J G 0.83fF
C5 En D 0.05fF
C6 Vref H 0.12fF
C7 w_16722_12162# C 0.12fF
C8 Vref A 0.81fF
C9 li_16144_1712# I 0.72fF
C10 li_16144_1712# En 0.05fF
C11 H w_16722_12162# 0.05fF
C12 w_16722_12162# A 0.03fF
C13 J En 0.47fF
C14 En A 0.42fF
C15 H C 0.06fF
C16 En G 0.39fF
C17 A C 0.66fF
C18 li_16144_1712# GND 3.98fF
C19 D GND 0.12fF
C20 B GND 0.69fF
C21 En GND 6.61fF
C22 C GND 5.08fF
C23 w_16722_12162# GND 59.23fF
C24 I GND 4.44fF
.ends
