magic
tech sky130A
magscale 1 2
timestamp 1620723023
<< nwell >>
rect 16722 12162 22724 13294
<< poly >>
rect 17212 7836 17562 7840
rect 17212 7790 22150 7836
rect 17212 7785 20645 7790
rect 17212 7683 17304 7785
rect 17406 7688 20645 7785
rect 20747 7688 22150 7790
rect 17406 7683 22150 7688
rect 17212 7652 22150 7683
rect 17212 7650 17566 7652
rect 18240 7650 18450 7652
rect 17212 7642 17562 7650
rect 20094 7644 20464 7652
rect 19492 6632 19828 6634
rect 18178 6630 19150 6632
rect 19370 6630 20754 6632
rect 18178 6545 20754 6630
rect 14302 6493 14504 6526
rect 14302 6459 14444 6493
rect 14478 6459 14504 6493
rect 14302 6432 14504 6459
rect 18178 6443 18755 6545
rect 18857 6443 20754 6545
rect 18178 6426 20754 6443
rect 18178 6346 19076 6426
rect 19136 6422 20754 6426
rect 19136 6418 19504 6422
rect 19812 6346 20754 6422
rect 14940 2342 15850 2390
rect 14940 2209 15846 2342
rect 14940 2107 15542 2209
rect 15644 2107 15846 2209
rect 14940 1992 15846 2107
rect 15294 1990 15846 1992
rect 16466 2144 17442 2422
rect 16466 2140 17864 2144
rect 21476 2140 22444 2308
rect 23092 2140 24068 2408
rect 24828 2366 25764 2374
rect 24828 2140 25784 2366
rect 16466 2017 25784 2140
rect 16466 1915 19161 2017
rect 19263 1915 25784 2017
rect 16466 1838 25784 1915
rect 16466 1836 24234 1838
rect 24828 1836 25784 1838
rect 16466 1826 17864 1836
<< polycont >>
rect 17304 7683 17406 7785
rect 20645 7688 20747 7790
rect 14444 6459 14478 6493
rect 18755 6443 18857 6545
rect 15542 2107 15644 2209
rect 19161 1915 19263 2017
<< locali >>
rect 16858 13121 17326 13124
rect 16858 13087 16861 13121
rect 16895 13087 16993 13121
rect 17027 13087 17149 13121
rect 17183 13087 17289 13121
rect 17323 13087 17326 13121
rect 16858 13086 17326 13087
rect 18920 13121 19372 13124
rect 18920 13087 18921 13121
rect 18955 13087 19069 13121
rect 19103 13087 19221 13121
rect 19255 13087 19337 13121
rect 19371 13087 19372 13121
rect 18920 13086 19372 13087
rect 20940 13121 21330 13124
rect 20940 13087 20943 13121
rect 20977 13087 21063 13121
rect 21097 13087 21189 13121
rect 21223 13087 21295 13121
rect 21329 13087 21330 13121
rect 20940 13086 21330 13087
rect 26730 13121 27246 13122
rect 26730 13087 26733 13121
rect 26767 13087 26903 13121
rect 26937 13087 27049 13121
rect 27083 13087 27211 13121
rect 27245 13087 27246 13121
rect 26730 13086 27246 13087
rect 17032 11698 17200 13086
rect 19034 11698 19202 13086
rect 21042 11690 21210 13086
rect 26866 11208 27030 13086
rect 26864 10462 27030 11208
rect 26864 10450 27010 10462
rect 2568 8616 3528 8742
rect 12242 8620 15822 8730
rect 2576 4330 2676 8616
rect 15702 8226 15818 8620
rect 15702 8208 15824 8226
rect 15712 7574 15824 8208
rect 17240 7785 17464 7826
rect 17240 7683 17304 7785
rect 17406 7683 17464 7785
rect 15632 7419 15970 7574
rect 15632 7313 15734 7419
rect 15840 7313 15970 7419
rect 15632 7158 15970 7313
rect 17240 7046 17464 7683
rect 18254 7222 18398 8176
rect 22240 8164 23056 8170
rect 20240 7340 20402 8020
rect 22240 7998 23062 8164
rect 20620 7790 20782 7836
rect 20620 7688 20645 7790
rect 20747 7688 20782 7790
rect 20620 7350 20782 7688
rect 20620 7340 20788 7350
rect 19580 7262 20788 7340
rect 16088 7044 17464 7046
rect 15920 7042 17464 7044
rect 18252 7110 19328 7222
rect 19568 7154 20788 7262
rect 19568 7148 20760 7154
rect 14386 6843 14530 6892
rect 14386 6809 14442 6843
rect 14476 6809 14530 6843
rect 14386 6756 14530 6809
rect 15920 6870 17460 7042
rect 18252 7040 19332 7110
rect 17882 6878 18096 6946
rect 18254 6878 18388 7040
rect 14426 6493 14500 6756
rect 14426 6459 14444 6493
rect 14478 6459 14500 6493
rect 14426 6432 14500 6459
rect 15920 6100 16088 6870
rect 17882 6858 18388 6878
rect 17882 6824 17963 6858
rect 17997 6850 18388 6858
rect 17997 6824 18382 6850
rect 17882 6786 18382 6824
rect 17882 6752 17963 6786
rect 17997 6752 18382 6786
rect 17882 6738 18382 6752
rect 17882 6676 18096 6738
rect 18704 6545 18896 7040
rect 18704 6443 18755 6545
rect 18857 6443 18896 6545
rect 18704 6398 18896 6443
rect 17532 6070 18014 6244
rect 19170 6170 19332 7040
rect 19568 6788 19760 7148
rect 19570 6172 19752 6788
rect 20836 6064 21374 6232
rect 22900 6062 23062 7998
rect 24066 7292 24388 7554
rect 24066 7258 24189 7292
rect 24223 7258 24388 7292
rect 24066 7220 24388 7258
rect 24066 7186 24189 7220
rect 24223 7186 24388 7220
rect 24066 6986 24388 7186
rect 24118 6154 24262 6986
rect 2532 4272 2700 4330
rect 2532 4238 2586 4272
rect 2620 4238 2700 4272
rect 2532 4192 2700 4238
rect 2550 3378 2650 3512
rect 3524 3378 3624 3512
rect 4582 3350 4682 3484
rect 5544 3358 5644 3492
rect 6578 3362 6674 3486
rect 5790 3328 6972 3334
rect 2214 3304 6972 3328
rect 1082 3298 6972 3304
rect 868 3290 6972 3298
rect 810 3004 6972 3290
rect 810 2984 1184 3004
rect 2214 3000 6972 3004
rect 810 568 1114 2984
rect 2536 2852 2636 2986
rect 3574 2868 3674 3000
rect 4590 2852 4690 2986
rect 5566 2864 5666 2998
rect 5790 2968 6972 3000
rect 6578 2870 6674 2968
rect 9610 2956 10054 2992
rect 9610 2922 9753 2956
rect 9787 2922 9825 2956
rect 9859 2922 9897 2956
rect 9931 2922 10054 2956
rect 9610 2880 10054 2922
rect 11040 2874 12092 3002
rect 11836 2810 12086 2874
rect 11152 1405 11256 1422
rect 11152 1371 11187 1405
rect 11221 1371 11256 1405
rect 11152 1333 11256 1371
rect 11152 1299 11187 1333
rect 11221 1299 11256 1333
rect 11152 1282 11256 1299
rect 11836 1072 12092 2810
rect 26866 2798 27014 3542
rect 26870 2754 27002 2798
rect 26874 2638 27002 2754
rect 13294 1072 13756 1206
rect 14222 1188 14280 2398
rect 14514 1838 14570 2404
rect 14452 1769 14606 1838
rect 14452 1735 14511 1769
rect 14545 1735 14606 1769
rect 14452 1656 14606 1735
rect 11824 1007 13756 1072
rect 11824 829 13431 1007
rect 13537 829 13756 1007
rect 11824 800 13756 829
rect 13294 690 13756 800
rect 14224 718 14280 1188
rect 14708 1492 14884 2576
rect 15494 2209 15700 2268
rect 15494 2107 15542 2209
rect 15644 2107 15700 2209
rect 15158 1802 15292 1864
rect 15494 1802 15700 2107
rect 16298 1944 16408 2528
rect 19076 2017 19334 2070
rect 15158 1765 15700 1802
rect 15158 1731 15197 1765
rect 15231 1731 15700 1765
rect 15158 1704 15700 1731
rect 16144 1831 16428 1944
rect 19076 1915 19161 2017
rect 19263 1915 19334 2017
rect 19076 1858 19334 1915
rect 22510 1890 22606 2540
rect 16144 1797 16262 1831
rect 16296 1797 16428 1831
rect 16144 1712 16428 1797
rect 22458 1802 22656 1890
rect 22458 1768 22550 1802
rect 22584 1768 22656 1802
rect 15158 1654 15292 1704
rect 15494 1612 15700 1704
rect 22458 1692 22656 1768
rect 24618 1626 24764 2636
rect 25854 2476 27006 2638
rect 21954 1612 24764 1626
rect 14224 670 14286 718
rect 804 66 1116 568
rect 14230 66 14286 670
rect 14708 612 14888 1492
rect 15494 1466 24764 1612
rect 15494 1464 16404 1466
rect 16492 1464 24764 1466
rect 15494 1454 15700 1464
rect 15840 1456 16404 1464
rect 21858 1454 24764 1464
rect 15002 1072 15288 1176
rect 19566 1076 19754 1082
rect 22352 1076 22706 1116
rect 19476 1074 22706 1076
rect 16918 1072 22706 1074
rect 15002 1011 22706 1072
rect 15002 976 22468 1011
rect 15002 942 15131 976
rect 15165 942 22468 976
rect 15002 905 22468 942
rect 22574 905 22706 1011
rect 15002 904 22706 905
rect 15002 870 15131 904
rect 15165 870 22706 904
rect 15002 844 22706 870
rect 15002 842 22390 844
rect 15002 728 15288 842
rect 16918 840 19796 842
rect 19476 836 19796 840
rect 14710 66 14882 612
rect 670 65 1246 66
rect 670 31 671 65
rect 705 31 761 65
rect 795 31 851 65
rect 885 31 941 65
rect 975 31 1031 65
rect 1065 31 1121 65
rect 1155 31 1211 65
rect 1245 31 1246 65
rect 670 30 1246 31
rect 14016 65 14532 66
rect 14016 31 14141 65
rect 14175 31 14231 65
rect 14265 31 14321 65
rect 14355 31 14532 65
rect 14016 30 14532 31
rect 14566 65 15070 66
rect 14566 31 14682 65
rect 14716 31 14771 65
rect 14805 31 14860 65
rect 14894 31 15070 65
rect 14566 30 15070 31
rect 15166 30 15672 66
rect 15714 30 16220 66
rect 16316 30 26422 66
<< viali >>
rect 16861 13087 16895 13121
rect 16993 13087 17027 13121
rect 17149 13087 17183 13121
rect 17289 13087 17323 13121
rect 18921 13087 18955 13121
rect 19069 13087 19103 13121
rect 19221 13087 19255 13121
rect 19337 13087 19371 13121
rect 20943 13087 20977 13121
rect 21063 13087 21097 13121
rect 21189 13087 21223 13121
rect 21295 13087 21329 13121
rect 26733 13087 26767 13121
rect 26903 13087 26937 13121
rect 27049 13087 27083 13121
rect 27211 13087 27245 13121
rect 15734 7313 15840 7419
rect 14442 6809 14476 6843
rect 17963 6824 17997 6858
rect 17963 6752 17997 6786
rect 24189 7258 24223 7292
rect 24189 7186 24223 7220
rect 2586 4238 2620 4272
rect 9753 2922 9787 2956
rect 9825 2922 9859 2956
rect 9897 2922 9931 2956
rect 11187 1371 11221 1405
rect 11187 1299 11221 1333
rect 14511 1735 14545 1769
rect 13431 829 13537 1007
rect 15197 1731 15231 1765
rect 16262 1797 16296 1831
rect 22550 1768 22584 1802
rect 15131 942 15165 976
rect 22468 905 22574 1011
rect 15131 870 15165 904
rect 671 31 705 65
rect 761 31 795 65
rect 851 31 885 65
rect 941 31 975 65
rect 1031 31 1065 65
rect 1121 31 1155 65
rect 1211 31 1245 65
rect 14141 31 14175 65
rect 14231 31 14265 65
rect 14321 31 14355 65
rect 14682 31 14716 65
rect 14771 31 14805 65
rect 14860 31 14894 65
<< metal1 >>
rect 0 13121 28540 13152
rect 0 13087 16861 13121
rect 16895 13087 16993 13121
rect 17027 13087 17149 13121
rect 17183 13087 17289 13121
rect 17323 13087 18921 13121
rect 18955 13087 19069 13121
rect 19103 13087 19221 13121
rect 19255 13087 19337 13121
rect 19371 13087 20943 13121
rect 20977 13087 21063 13121
rect 21097 13087 21189 13121
rect 21223 13087 21295 13121
rect 21329 13087 26733 13121
rect 26767 13087 26903 13121
rect 26937 13087 27049 13121
rect 27083 13087 27211 13121
rect 27245 13087 28540 13121
rect 0 13056 28540 13087
rect 15632 7424 15970 7574
rect 15632 7419 15761 7424
rect 15813 7419 15970 7424
rect 15632 7313 15734 7419
rect 15840 7313 15970 7419
rect 15632 7308 15761 7313
rect 15813 7308 15970 7313
rect 15632 7158 15970 7308
rect 24066 7292 24388 7554
rect 24066 7265 24189 7292
rect 24223 7265 24388 7292
rect 24066 7213 24180 7265
rect 24232 7213 24388 7265
rect 24066 7186 24189 7213
rect 24223 7186 24388 7213
rect 24066 6986 24388 7186
rect 14386 6852 14530 6892
rect 14386 6800 14433 6852
rect 14485 6800 14530 6852
rect 14386 6756 14530 6800
rect 17882 6863 18096 6946
rect 17882 6811 17954 6863
rect 18006 6811 18096 6863
rect 17882 6799 18096 6811
rect 17882 6747 17954 6799
rect 18006 6747 18096 6799
rect 17882 6676 18096 6747
rect 2532 4272 2700 4330
rect 2532 4238 2586 4272
rect 2620 4238 2700 4272
rect 2532 4192 2700 4238
rect 2554 3668 2656 4192
rect 6564 3732 9810 3736
rect 3516 3638 9810 3732
rect 3568 2732 3646 3638
rect 6564 3608 9810 3638
rect 9388 3600 9810 3608
rect 9654 3012 9810 3600
rect 9654 2992 10016 3012
rect 9610 2956 10054 2992
rect 9610 2922 9753 2956
rect 9787 2922 9825 2956
rect 9859 2922 9897 2956
rect 9931 2922 10054 2956
rect 9610 2880 10054 2922
rect 2518 2638 5568 2732
rect 6554 2636 9142 2758
rect 9046 1396 9136 2636
rect 14454 1836 14514 1840
rect 14570 1836 14606 1840
rect 14454 1774 14606 1836
rect 14454 1722 14504 1774
rect 14556 1722 14606 1774
rect 14454 1656 14606 1722
rect 15154 1824 15294 1864
rect 16144 1840 16428 1944
rect 15154 1773 15298 1824
rect 15154 1721 15197 1773
rect 15249 1721 15298 1773
rect 15154 1708 15298 1721
rect 16144 1788 16253 1840
rect 16305 1788 16428 1840
rect 16144 1712 16428 1788
rect 22458 1886 22510 1888
rect 22606 1886 22658 1888
rect 22458 1812 22658 1886
rect 22458 1760 22542 1812
rect 22594 1760 22658 1812
rect 15154 1652 15294 1708
rect 22458 1688 22658 1760
rect 11038 1405 11398 1608
rect 11038 1396 11187 1405
rect 9046 1371 11187 1396
rect 11221 1371 11398 1405
rect 9046 1333 11398 1371
rect 9046 1299 11187 1333
rect 11221 1299 11398 1333
rect 9046 1262 11398 1299
rect 9052 1256 11398 1262
rect 11038 1120 11398 1256
rect 13300 1036 13758 1206
rect 13292 1007 13758 1036
rect 13292 832 13429 1007
rect 13300 827 13429 832
rect 13545 827 13758 1007
rect 13300 690 13758 827
rect 15004 1068 15292 1170
rect 22352 1068 22706 1116
rect 15004 982 15294 1068
rect 15004 930 15130 982
rect 15182 930 15294 982
rect 15004 918 15294 930
rect 15004 866 15130 918
rect 15182 866 15294 918
rect 15004 848 15294 866
rect 22350 1011 22706 1068
rect 22350 905 22468 1011
rect 22574 905 22706 1011
rect 22350 848 22706 905
rect 15004 728 15292 848
rect 22352 844 22706 848
rect 0 65 28540 96
rect 0 31 671 65
rect 705 31 761 65
rect 795 31 851 65
rect 885 31 941 65
rect 975 31 1031 65
rect 1065 31 1121 65
rect 1155 31 1211 65
rect 1245 31 14141 65
rect 14175 31 14231 65
rect 14265 31 14321 65
rect 14355 31 14682 65
rect 14716 31 14771 65
rect 14805 31 14860 65
rect 14894 31 28540 65
rect 0 0 28540 31
<< via1 >>
rect 15761 7419 15813 7424
rect 15761 7372 15813 7419
rect 15761 7313 15813 7360
rect 15761 7308 15813 7313
rect 24180 7258 24189 7265
rect 24189 7258 24223 7265
rect 24223 7258 24232 7265
rect 24180 7220 24232 7258
rect 24180 7213 24189 7220
rect 24189 7213 24223 7220
rect 24223 7213 24232 7220
rect 14433 6843 14485 6852
rect 14433 6809 14442 6843
rect 14442 6809 14476 6843
rect 14476 6809 14485 6843
rect 14433 6800 14485 6809
rect 17954 6858 18006 6863
rect 17954 6824 17963 6858
rect 17963 6824 17997 6858
rect 17997 6824 18006 6858
rect 17954 6811 18006 6824
rect 17954 6786 18006 6799
rect 17954 6752 17963 6786
rect 17963 6752 17997 6786
rect 17997 6752 18006 6786
rect 17954 6747 18006 6752
rect 14504 1769 14556 1774
rect 14504 1735 14511 1769
rect 14511 1735 14545 1769
rect 14545 1735 14556 1769
rect 14504 1722 14556 1735
rect 15197 1765 15249 1773
rect 15197 1731 15231 1765
rect 15231 1731 15249 1765
rect 15197 1721 15249 1731
rect 16253 1831 16305 1840
rect 16253 1797 16262 1831
rect 16262 1797 16296 1831
rect 16296 1797 16305 1831
rect 16253 1788 16305 1797
rect 22542 1802 22594 1812
rect 22542 1768 22550 1802
rect 22550 1768 22584 1802
rect 22584 1768 22594 1802
rect 22542 1760 22594 1768
rect 13429 829 13431 1007
rect 13431 829 13537 1007
rect 13537 829 13545 1007
rect 13429 827 13545 829
rect 15130 976 15182 982
rect 15130 942 15131 976
rect 15131 942 15165 976
rect 15165 942 15182 976
rect 15130 930 15182 942
rect 15130 904 15182 918
rect 15130 870 15131 904
rect 15131 870 15165 904
rect 15165 870 15182 904
rect 15130 866 15182 870
rect 22495 931 22547 983
<< metal2 >>
rect 15632 7424 15970 7574
rect 15632 7372 15761 7424
rect 15813 7372 15970 7424
rect 15632 7360 15970 7372
rect 15632 7308 15761 7360
rect 15813 7334 15970 7360
rect 24066 7334 24388 7554
rect 15813 7308 24388 7334
rect 15632 7265 24388 7308
rect 15632 7213 24180 7265
rect 24232 7213 24388 7265
rect 15632 7204 24388 7213
rect 15632 7158 15970 7204
rect 24066 6986 24388 7204
rect 14386 6852 14530 6892
rect 14386 6800 14433 6852
rect 14485 6844 14530 6852
rect 17882 6863 18096 6946
rect 17882 6844 17954 6863
rect 14485 6811 17954 6844
rect 18006 6811 18096 6863
rect 14485 6800 18096 6811
rect 14386 6799 18096 6800
rect 14386 6790 17954 6799
rect 14386 6756 14530 6790
rect 15902 6786 16130 6790
rect 17882 6747 17954 6790
rect 18006 6747 18096 6799
rect 17882 6676 18096 6747
rect 14454 1836 14514 1840
rect 14570 1836 14606 1840
rect 14454 1820 14606 1836
rect 15154 1820 15294 1864
rect 14454 1774 15294 1820
rect 14454 1722 14504 1774
rect 14556 1773 15294 1774
rect 14556 1722 15197 1773
rect 14454 1721 15197 1722
rect 15249 1721 15294 1773
rect 14454 1692 15294 1721
rect 16144 1840 16428 1944
rect 16144 1788 16253 1840
rect 16305 1788 16428 1840
rect 16144 1712 16428 1788
rect 22458 1886 22510 1888
rect 22606 1886 22658 1888
rect 22458 1812 22658 1886
rect 22458 1760 22542 1812
rect 22594 1760 22658 1812
rect 14454 1656 14606 1692
rect 14692 1690 14948 1692
rect 15154 1652 15294 1692
rect 11038 1410 11398 1608
rect 16234 1410 16382 1712
rect 22458 1688 22658 1760
rect 11038 1270 16386 1410
rect 22494 1320 22572 1688
rect 11038 1120 11398 1270
rect 16234 1262 16382 1270
rect 13300 1084 13758 1206
rect 14214 1084 14318 1086
rect 15004 1084 15292 1170
rect 22496 1116 22572 1320
rect 13300 1007 15292 1084
rect 13300 827 13429 1007
rect 13545 982 15292 1007
rect 13545 930 15130 982
rect 15182 930 15292 982
rect 13545 918 15292 930
rect 13545 866 15130 918
rect 15182 866 15292 918
rect 13545 827 15292 866
rect 22352 983 22706 1116
rect 22352 931 22495 983
rect 22547 931 22706 983
rect 22352 844 22706 931
rect 13300 796 15292 827
rect 13300 690 13758 796
rect 15004 728 15292 796
use resistor30K  resistor30K_0
timestamp 1620719712
transform 1 0 10016 0 1 2900
box -402 -22 1462 96
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_5
timestamp 1615375237
transform 1 0 6218 0 1 2296
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_6
timestamp 1615375237
transform 1 0 5200 0 1 2284
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_7
timestamp 1615375237
transform 1 0 4230 0 1 2284
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_8
timestamp 1615375237
transform 1 0 3226 0 1 2296
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_9
timestamp 1615375237
transform 1 0 2182 0 1 2266
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_3
timestamp 1615375237
transform 1 0 3180 0 1 3292
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_4
timestamp 1615375237
transform 1 0 2206 0 1 3292
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_0
timestamp 1615375237
transform 1 0 6218 0 1 3270
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_1
timestamp 1615375237
transform 1 0 5198 0 1 3270
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_2
timestamp 1615375237
transform 1 0 4224 0 1 3270
box 26 26 770 795
use resistor273K  resistor273K_0
timestamp 1620719712
transform 1 0 3522 0 1 8642
box -430 -10 9170 80
use nmos2metal120  nmos2metal120_1
timestamp 1620722909
transform 1 0 14524 0 1 2410
box -16 -16 50 50
use nmos2metal120  nmos2metal120_0
timestamp 1620722909
transform 1 0 14238 0 1 2406
box -16 -16 50 50
use nmos_substrate  nmos_substrate_21
timestamp 1620719712
transform 1 0 14470 0 1 0
box -26 -26 122 122
use nmos_substrate  nmos_substrate_20
timestamp 1620719712
transform 1 0 13920 0 1 0
box -26 -26 122 122
use nmos_substrate  nmos_substrate_19
timestamp 1620719712
transform 1 0 15070 0 1 0
box -26 -26 122 122
use nmos_substrate  nmos_substrate_18
timestamp 1620719712
transform 1 0 15620 0 1 0
box -26 -26 122 122
use NMOS520  NMOS520_6
timestamp 1620719712
transform 1 0 14910 0 1 2360
box -202 -100 1202 4100
use NMOS120  NMOS120_0
timestamp 1620719712
transform 1 0 14302 0 1 2380
box -80 -60 280 4060
use nmos2metal  nmos2metal_13
timestamp 1620719712
transform 1 0 14708 0 1 2456
box 0 0 200 200
use nmos_substrate  nmos_substrate_17
timestamp 1620719712
transform 1 0 16220 0 1 0
box -26 -26 122 122
use nmos_substrate  nmos_substrate_16
timestamp 1620719712
transform 1 0 16820 0 1 0
box -26 -26 122 122
use nmos_substrate  nmos_substrate_15
timestamp 1620719712
transform 1 0 17420 0 1 0
box -26 -26 122 122
use NMOS520  NMOS520_5
timestamp 1620719712
transform 1 0 16458 0 1 2350
box -202 -100 1202 4100
use nmos2metal  nmos2metal_12
timestamp 1620719712
transform 1 0 16260 0 1 2454
box 0 0 200 200
use nmos_substrate  nmos_substrate_14
timestamp 1620719712
transform 1 0 19220 0 1 0
box -26 -26 122 122
use nmos_substrate  nmos_substrate_13
timestamp 1620719712
transform 1 0 18620 0 1 0
box -26 -26 122 122
use nmos_substrate  nmos_substrate_12
timestamp 1620719712
transform 1 0 18020 0 1 0
box -26 -26 122 122
use nmos_substrate  nmos_substrate_11
timestamp 1620719712
transform 1 0 19820 0 1 0
box -26 -26 122 122
use NMOS520  NMOS520_3
timestamp 1620719712
transform 1 0 18150 0 1 2350
box -202 -100 1202 4100
use NMOS520  NMOS520_4
timestamp 1620719712
transform 1 0 19758 0 1 2350
box -202 -100 1202 4100
use nmos_substrate  nmos_substrate_10
timestamp 1620719712
transform 1 0 21020 0 1 0
box -26 -26 122 122
use nmos_substrate  nmos_substrate_9
timestamp 1620719712
transform 1 0 20420 0 1 0
box -26 -26 122 122
use NMOS520  NMOS520_2
timestamp 1620719712
transform 1 0 21446 0 1 2360
box -202 -100 1202 4100
use PMOS520  PMOS520_2
timestamp 1620719712
transform 1 0 17220 0 1 7896
box -502 -372 1500 4374
use nmos2metal  nmos2metal_10
timestamp 1620719712
transform 1 0 15906 0 1 6062
box 0 0 200 200
use nmos2metal  nmos2metal_11
timestamp 1620719712
transform 1 0 17462 0 1 6056
box 0 0 200 200
use pmos2metaal  pmos2metaal_5
timestamp 1620719712
transform 1 0 18224 0 1 8002
box -72 -66 272 268
use PMOS520  PMOS520_1
timestamp 1620719712
transform 1 0 19218 0 1 7886
box -502 -372 1500 4374
use nmos2metal  nmos2metal_7
timestamp 1620719712
transform 1 0 17948 0 1 6054
box 0 0 200 200
use nmos2metal  nmos2metal_8
timestamp 1620719712
transform 1 0 19558 0 1 6054
box 0 0 200 200
use nmos2metal  nmos2metal_9
timestamp 1620719712
transform 1 0 19148 0 1 6054
box 0 0 200 200
use pmos2metaal  pmos2metaal_4
timestamp 1620719712
transform 1 0 20216 0 1 7982
box -72 -66 272 268
use PMOS520  PMOS520_0
timestamp 1620719712
transform 1 0 21214 0 1 7884
box -502 -372 1500 4374
use nmos2metal  nmos2metal_5
timestamp 1620719712
transform 1 0 21248 0 1 6054
box 0 0 200 200
use nmos2metal  nmos2metal_6
timestamp 1620719712
transform 1 0 20760 0 1 6046
box 0 0 200 200
use pmos2metaal  pmos2metaal_3
timestamp 1620719712
transform 1 0 17014 0 1 11590
box -72 -66 272 268
use pmos_substrate  pmos_substrate_5
timestamp 1620719712
transform 1 0 17606 0 1 13056
box -66 -68 162 162
use pmos2metaal  pmos2metaal_2
timestamp 1620719712
transform 1 0 19014 0 1 11582
box -72 -66 272 268
use pmos_substrate  pmos_substrate_4
timestamp 1620719712
transform 1 0 19656 0 1 13056
box -66 -68 162 162
use pmos_substrate  pmos_substrate_3
timestamp 1620719712
transform 1 0 18290 0 1 13056
box -66 -68 162 162
use pmos2metaal  pmos2metaal_1
timestamp 1620719712
transform 1 0 21014 0 1 11580
box -72 -66 272 268
use pmos_substrate  pmos_substrate_2
timestamp 1620719712
transform 1 0 20226 0 1 13056
box -66 -68 162 162
use pmos2metaal  pmos2metaal_0
timestamp 1620719712
transform 1 0 22206 0 1 7980
box -72 -66 272 268
use nmos_substrate  nmos_substrate_8
timestamp 1620719712
transform 1 0 22218 0 1 0
box -26 -26 122 122
use nmos_substrate  nmos_substrate_7
timestamp 1620719712
transform 1 0 21620 0 1 0
box -26 -26 122 122
use pmos_substrate  pmos_substrate_1
timestamp 1620719712
transform 1 0 22062 0 1 13056
box -66 -68 162 162
use pmos_substrate  pmos_substrate_0
timestamp 1620719712
transform 1 0 21496 0 1 13056
box -66 -68 162 162
use nmos_substrate  nmos_substrate_6
timestamp 1620719712
transform 1 0 22820 0 1 0
box -26 -26 122 122
use nmos2metal  nmos2metal_4
timestamp 1620719712
transform 1 0 22454 0 1 2462
box 0 0 200 200
use nmos_substrate  nmos_substrate_5
timestamp 1620719712
transform 1 0 23420 0 1 0
box -26 -26 122 122
use nmos_substrate  nmos_substrate_4
timestamp 1620719712
transform 1 0 24020 0 1 0
box -26 -26 122 122
use NMOS520  NMOS520_1
timestamp 1620719712
transform 1 0 23088 0 1 2350
box -202 -100 1202 4100
use nmos2metal  nmos2metal_2
timestamp 1620719712
transform 1 0 22882 0 1 6034
box 0 0 200 200
use nmos2metal  nmos2metal_3
timestamp 1620719712
transform 1 0 24092 0 1 6026
box 0 0 200 200
use nmos_substrate  nmos_substrate_3
timestamp 1620719712
transform 1 0 25220 0 1 0
box -26 -26 122 122
use nmos_substrate  nmos_substrate_2
timestamp 1620719712
transform 1 0 24620 0 1 0
box -26 -26 122 122
use NMOS520  NMOS520_0
timestamp 1620719712
transform 1 0 24788 0 1 2360
box -202 -100 1202 4100
use nmos2metal  nmos2metal_1
timestamp 1620719712
transform 1 0 24592 0 1 2460
box 0 0 200 200
use resistor200K  resistor200K_0
timestamp 1620719712
transform 0 1 26910 -1 0 10506
box -700 -40 7704 102
use nmos_substrate  nmos_substrate_1
timestamp 1620719712
transform 1 0 25820 0 1 0
box -26 -26 122 122
use nmos_substrate  nmos_substrate_0
timestamp 1620719712
transform 1 0 26420 0 1 0
box -26 -26 122 122
use nmos2metal  nmos2metal_0
timestamp 1620719712
transform 1 0 25790 0 1 2458
box 0 0 200 200
<< labels >>
flabel poly s 19936 6370 20158 6624 0 FreeSans 3125 0 0 0 A
flabel metal1 s 8076 3704 8076 3704 0 FreeSans 3125 0 0 0 E
rlabel poly s 21236 7726 21236 7726 4 C
flabel locali s 22970 7622 22970 7622 0 FreeSans 3125 0 0 0 H
rlabel poly s 20276 6456 20276 6456 4 A
rlabel poly s 18652 7708 18652 7708 4 C
rlabel locali s 17818 6132 17818 6132 4 B
rlabel locali s 21130 6132 21130 6132 4 D
rlabel locali s 11914 2476 11914 2476 4 J
rlabel metal1 s 8714 3658 8714 3658 4 E
rlabel metal1 s 8372 2686 8372 2686 4 I
rlabel locali s 26510 2526 26510 2526 4 K
rlabel locali s 21532 1524 21532 1524 4 G
rlabel locali s 2630 5638 2630 5638 4 F
flabel metal1 s 11202 36 11202 36 0 FreeSans 3125 0 0 0 GND
port 1 nsew
flabel locali s 13292 8670 13292 8670 0 FreeSans 3125 0 0 0 Vref
port 2 nsew
flabel locali s 19130 1888 19294 2044 0 FreeSans 3125 0 0 0 En
port 3 nsew
flabel metal1 s 9822 13102 9822 13102 0 FreeSans 2000 0 0 0 VDD
port 4 nsew
<< properties >>
string FIXED_BBOX 0 48 28540 13104
<< end >>
