magic
tech sky130A
timestamp 1619503262
<< error_p >>
rect 84 94 90 96
rect 6 90 94 94
rect 4 86 96 90
rect 4 84 14 86
rect 10 14 14 84
rect 86 84 96 86
rect 86 14 94 84
rect 10 10 94 14
rect 84 6 94 10
rect 84 4 90 6
<< mvndiffc >>
rect 10 10 90 90
<< locali >>
rect 0 90 100 100
rect 0 10 10 90
rect 90 10 100 90
rect 0 0 100 10
<< end >>
