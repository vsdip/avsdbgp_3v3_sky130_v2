magic
tech sky130A
timestamp 1615565174
<< mvnmos >>
rect 1100 0 1600 2000
<< mvndiff >>
rect 1000 0 1100 2000
rect 1600 0 1700 2000
<< poly >>
rect 1100 2000 1600 2050
rect 1100 -50 1600 0
<< end >>
