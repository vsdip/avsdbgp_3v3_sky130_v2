VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO BGR
  CLASS BLOCK ;
  FOREIGN BGR ;
  ORIGIN 0.000 -0.240 ;
  SIZE 142.700 BY 65.280 ;
  PIN GND
    ANTENNAGATEAREA 60.024998 ;
    ANTENNADIFFAREA 122.928795 ;
    PORT
      LAYER pwell ;
        RECT 11.160 19.805 14.880 20.310 ;
        RECT 11.160 17.095 11.665 19.805 ;
        RECT 14.375 17.095 14.880 19.805 ;
        RECT 11.160 16.590 14.880 17.095 ;
        RECT 16.030 19.805 19.750 20.310 ;
        RECT 16.030 17.095 16.535 19.805 ;
        RECT 19.245 17.095 19.750 19.805 ;
        RECT 16.030 16.590 19.750 17.095 ;
        RECT 21.250 19.695 24.970 20.200 ;
        RECT 21.250 16.985 21.755 19.695 ;
        RECT 24.465 16.985 24.970 19.695 ;
        RECT 21.250 16.480 24.970 16.985 ;
        RECT 26.120 19.695 29.840 20.200 ;
        RECT 26.120 16.985 26.625 19.695 ;
        RECT 29.335 16.985 29.840 19.695 ;
        RECT 26.120 16.480 29.840 16.985 ;
        RECT 31.220 19.695 34.940 20.200 ;
        RECT 31.220 16.985 31.725 19.695 ;
        RECT 34.435 16.985 34.940 19.695 ;
        RECT 31.220 16.480 34.940 16.985 ;
        RECT 11.040 14.675 14.760 15.180 ;
        RECT 11.040 11.965 11.545 14.675 ;
        RECT 14.255 11.965 14.760 14.675 ;
        RECT 11.040 11.460 14.760 11.965 ;
        RECT 16.260 14.825 19.980 15.330 ;
        RECT 16.260 12.115 16.765 14.825 ;
        RECT 19.475 12.115 19.980 14.825 ;
        RECT 16.260 11.610 19.980 12.115 ;
        RECT 21.280 14.765 25.000 15.270 ;
        RECT 21.280 12.055 21.785 14.765 ;
        RECT 24.495 12.055 25.000 14.765 ;
        RECT 21.280 11.550 25.000 12.055 ;
        RECT 26.130 14.765 29.850 15.270 ;
        RECT 26.130 12.055 26.635 14.765 ;
        RECT 29.345 12.055 29.850 14.765 ;
        RECT 26.130 11.550 29.850 12.055 ;
        RECT 31.220 14.825 34.940 15.330 ;
        RECT 31.220 12.115 31.725 14.825 ;
        RECT 34.435 12.115 34.940 14.825 ;
        RECT 31.220 11.610 34.940 12.115 ;
        RECT 69.470 -0.130 70.210 0.610 ;
        RECT 72.220 -0.130 72.960 0.610 ;
        RECT 75.220 -0.130 75.960 0.610 ;
        RECT 77.970 -0.130 78.710 0.610 ;
        RECT 80.970 -0.130 81.710 0.610 ;
        RECT 83.970 -0.130 84.710 0.610 ;
        RECT 86.970 -0.130 87.710 0.610 ;
        RECT 89.970 -0.130 90.710 0.610 ;
        RECT 92.970 -0.130 93.710 0.610 ;
        RECT 95.970 -0.130 96.710 0.610 ;
        RECT 98.970 -0.130 99.710 0.610 ;
        RECT 101.970 -0.130 102.710 0.610 ;
        RECT 104.970 -0.130 105.710 0.610 ;
        RECT 107.970 -0.130 108.710 0.610 ;
        RECT 110.960 -0.130 111.700 0.610 ;
        RECT 113.970 -0.130 114.710 0.610 ;
        RECT 116.970 -0.130 117.710 0.610 ;
        RECT 119.970 -0.130 120.710 0.610 ;
        RECT 122.970 -0.130 123.710 0.610 ;
        RECT 125.970 -0.130 126.710 0.610 ;
        RECT 128.970 -0.130 129.710 0.610 ;
        RECT 131.970 -0.130 132.710 0.610 ;
      LAYER li1 ;
        RECT 11.160 19.805 14.880 20.310 ;
        RECT 11.160 17.095 11.665 19.805 ;
        RECT 11.975 19.135 14.065 19.495 ;
        RECT 11.975 17.765 12.335 19.135 ;
        RECT 13.705 17.765 14.065 19.135 ;
        RECT 11.975 17.405 14.065 17.765 ;
        RECT 12.750 17.095 13.250 17.405 ;
        RECT 14.375 17.095 14.880 19.805 ;
        RECT 11.160 16.640 14.880 17.095 ;
        RECT 16.030 19.805 19.750 20.310 ;
        RECT 16.030 17.095 16.535 19.805 ;
        RECT 16.845 19.135 18.935 19.495 ;
        RECT 16.845 17.765 17.205 19.135 ;
        RECT 18.575 17.765 18.935 19.135 ;
        RECT 16.845 17.405 18.935 17.765 ;
        RECT 17.620 17.095 18.120 17.405 ;
        RECT 19.245 17.095 19.750 19.805 ;
        RECT 16.030 16.640 19.750 17.095 ;
        RECT 21.250 19.695 24.970 20.200 ;
        RECT 21.250 16.985 21.755 19.695 ;
        RECT 22.065 19.025 24.155 19.385 ;
        RECT 22.065 17.655 22.425 19.025 ;
        RECT 23.795 17.655 24.155 19.025 ;
        RECT 22.065 17.295 24.155 17.655 ;
        RECT 22.910 16.985 23.410 17.295 ;
        RECT 24.465 16.985 24.970 19.695 ;
        RECT 21.250 16.640 24.970 16.985 ;
        RECT 26.120 19.695 29.840 20.200 ;
        RECT 26.120 16.985 26.625 19.695 ;
        RECT 26.935 19.025 29.025 19.385 ;
        RECT 26.935 17.655 27.295 19.025 ;
        RECT 28.665 17.655 29.025 19.025 ;
        RECT 26.935 17.295 29.025 17.655 ;
        RECT 27.720 16.985 28.220 17.295 ;
        RECT 29.335 16.985 29.840 19.695 ;
        RECT 26.120 16.670 29.840 16.985 ;
        RECT 31.220 19.695 34.940 20.200 ;
        RECT 31.220 16.985 31.725 19.695 ;
        RECT 32.035 19.025 34.125 19.385 ;
        RECT 32.035 17.655 32.395 19.025 ;
        RECT 33.765 17.655 34.125 19.025 ;
        RECT 32.035 17.295 34.125 17.655 ;
        RECT 32.890 16.985 33.370 17.295 ;
        RECT 34.435 16.985 34.940 19.695 ;
        RECT 31.220 16.670 34.940 16.985 ;
        RECT 26.120 16.640 34.940 16.670 ;
        RECT 11.070 16.520 34.940 16.640 ;
        RECT 5.410 16.490 34.940 16.520 ;
        RECT 4.340 16.480 34.940 16.490 ;
        RECT 4.340 16.450 34.860 16.480 ;
        RECT 4.050 15.330 34.860 16.450 ;
        RECT 4.050 15.020 34.940 15.330 ;
        RECT 4.050 14.920 5.920 15.020 ;
        RECT 11.040 15.000 34.940 15.020 ;
        RECT 4.050 2.840 5.570 14.920 ;
        RECT 11.040 14.675 14.760 15.000 ;
        RECT 11.040 11.965 11.545 14.675 ;
        RECT 12.680 14.365 13.180 14.675 ;
        RECT 11.855 14.005 13.945 14.365 ;
        RECT 11.855 12.635 12.215 14.005 ;
        RECT 13.585 12.635 13.945 14.005 ;
        RECT 11.855 12.275 13.945 12.635 ;
        RECT 14.255 11.965 14.760 14.675 ;
        RECT 11.040 11.460 14.760 11.965 ;
        RECT 16.260 14.825 19.980 15.000 ;
        RECT 16.260 12.115 16.765 14.825 ;
        RECT 17.870 14.515 18.370 14.825 ;
        RECT 17.075 14.155 19.165 14.515 ;
        RECT 17.075 12.785 17.435 14.155 ;
        RECT 18.805 12.785 19.165 14.155 ;
        RECT 17.075 12.425 19.165 12.785 ;
        RECT 19.475 12.115 19.980 14.825 ;
        RECT 16.260 11.610 19.980 12.115 ;
        RECT 21.280 14.765 25.000 15.000 ;
        RECT 21.280 12.055 21.785 14.765 ;
        RECT 22.950 14.455 23.450 14.765 ;
        RECT 22.095 14.095 24.185 14.455 ;
        RECT 22.095 12.725 22.455 14.095 ;
        RECT 23.825 12.725 24.185 14.095 ;
        RECT 22.095 12.365 24.185 12.725 ;
        RECT 24.495 12.055 25.000 14.765 ;
        RECT 21.280 11.550 25.000 12.055 ;
        RECT 26.130 14.840 34.940 15.000 ;
        RECT 26.130 14.765 29.850 14.840 ;
        RECT 26.130 12.055 26.635 14.765 ;
        RECT 27.830 14.455 28.330 14.765 ;
        RECT 26.945 14.095 29.035 14.455 ;
        RECT 26.945 12.725 27.305 14.095 ;
        RECT 28.675 12.725 29.035 14.095 ;
        RECT 26.945 12.365 29.035 12.725 ;
        RECT 29.345 12.055 29.850 14.765 ;
        RECT 26.130 11.550 29.850 12.055 ;
        RECT 31.220 14.825 34.940 14.840 ;
        RECT 31.220 12.115 31.725 14.825 ;
        RECT 32.890 14.515 33.370 14.825 ;
        RECT 32.035 14.155 34.125 14.515 ;
        RECT 32.035 12.785 32.395 14.155 ;
        RECT 33.765 12.785 34.125 14.155 ;
        RECT 32.035 12.425 34.125 12.785 ;
        RECT 34.435 12.115 34.940 14.825 ;
        RECT 73.540 12.280 74.540 13.280 ;
        RECT 31.220 11.610 34.940 12.115 ;
        RECT 71.110 11.950 71.440 12.280 ;
        RECT 71.110 5.940 71.400 11.950 ;
        RECT 71.120 3.590 71.400 5.940 ;
        RECT 73.540 7.460 74.420 12.280 ;
        RECT 71.120 3.350 71.430 3.590 ;
        RECT 4.020 0.330 5.580 2.840 ;
        RECT 69.600 0.330 70.080 0.480 ;
        RECT 71.150 0.330 71.430 3.350 ;
        RECT 73.540 3.060 74.440 7.460 ;
        RECT 72.350 0.330 72.830 0.480 ;
        RECT 73.550 0.330 74.410 3.060 ;
        RECT 75.350 0.330 75.830 0.480 ;
        RECT 78.100 0.330 78.580 0.480 ;
        RECT 81.100 0.330 81.580 0.480 ;
        RECT 84.100 0.330 84.580 0.480 ;
        RECT 87.100 0.330 87.580 0.480 ;
        RECT 90.100 0.330 90.580 0.480 ;
        RECT 93.100 0.330 93.580 0.480 ;
        RECT 96.100 0.330 96.580 0.480 ;
        RECT 99.100 0.330 99.580 0.480 ;
        RECT 102.100 0.330 102.580 0.480 ;
        RECT 105.100 0.330 105.580 0.480 ;
        RECT 108.100 0.330 108.580 0.480 ;
        RECT 111.090 0.330 111.570 0.480 ;
        RECT 114.100 0.330 114.580 0.480 ;
        RECT 117.100 0.330 117.580 0.480 ;
        RECT 120.100 0.330 120.580 0.480 ;
        RECT 123.100 0.330 123.580 0.480 ;
        RECT 126.100 0.330 126.580 0.480 ;
        RECT 129.100 0.330 129.580 0.480 ;
        RECT 132.100 0.330 132.580 0.480 ;
        RECT 3.350 0.150 6.230 0.330 ;
        RECT 69.600 0.150 132.580 0.330 ;
        RECT 69.600 0.000 70.080 0.150 ;
        RECT 72.350 0.000 72.830 0.150 ;
        RECT 75.350 0.000 75.830 0.150 ;
        RECT 78.100 0.000 78.580 0.150 ;
        RECT 81.100 0.000 81.580 0.150 ;
        RECT 84.100 0.000 84.580 0.150 ;
        RECT 87.100 0.000 87.580 0.150 ;
        RECT 90.100 0.000 90.580 0.150 ;
        RECT 93.100 0.000 93.580 0.150 ;
        RECT 96.100 0.000 96.580 0.150 ;
        RECT 99.100 0.000 99.580 0.150 ;
        RECT 102.100 0.000 102.580 0.150 ;
        RECT 105.100 0.000 105.580 0.150 ;
        RECT 108.100 0.000 108.580 0.150 ;
        RECT 111.090 0.000 111.570 0.150 ;
        RECT 114.100 0.000 114.580 0.150 ;
        RECT 117.100 0.000 117.580 0.150 ;
        RECT 120.100 0.000 120.580 0.150 ;
        RECT 123.100 0.000 123.580 0.150 ;
        RECT 126.100 0.000 126.580 0.150 ;
        RECT 129.100 0.000 129.580 0.150 ;
        RECT 132.100 0.000 132.580 0.150 ;
      LAYER mcon ;
        RECT 3.355 0.155 3.525 0.325 ;
        RECT 3.805 0.155 3.975 0.325 ;
        RECT 4.255 0.155 4.425 0.325 ;
        RECT 4.705 0.155 4.875 0.325 ;
        RECT 5.155 0.155 5.325 0.325 ;
        RECT 5.605 0.155 5.775 0.325 ;
        RECT 6.055 0.155 6.225 0.325 ;
        RECT 69.750 0.150 69.920 0.320 ;
        RECT 70.705 0.155 70.875 0.325 ;
        RECT 71.155 0.155 71.325 0.325 ;
        RECT 71.605 0.155 71.775 0.325 ;
        RECT 72.500 0.150 72.670 0.320 ;
        RECT 73.410 0.155 73.580 0.325 ;
        RECT 73.855 0.155 74.025 0.325 ;
        RECT 74.300 0.155 74.470 0.325 ;
        RECT 75.500 0.150 75.670 0.320 ;
        RECT 78.250 0.150 78.420 0.320 ;
        RECT 81.250 0.150 81.420 0.320 ;
        RECT 84.250 0.150 84.420 0.320 ;
        RECT 87.250 0.150 87.420 0.320 ;
        RECT 90.250 0.150 90.420 0.320 ;
        RECT 93.250 0.150 93.420 0.320 ;
        RECT 96.250 0.150 96.420 0.320 ;
        RECT 99.250 0.150 99.420 0.320 ;
        RECT 102.250 0.150 102.420 0.320 ;
        RECT 105.250 0.150 105.420 0.320 ;
        RECT 108.250 0.150 108.420 0.320 ;
        RECT 111.240 0.150 111.410 0.320 ;
        RECT 114.250 0.150 114.420 0.320 ;
        RECT 117.250 0.150 117.420 0.320 ;
        RECT 120.250 0.150 120.420 0.320 ;
        RECT 123.250 0.150 123.420 0.320 ;
        RECT 126.250 0.150 126.420 0.320 ;
        RECT 129.250 0.150 129.420 0.320 ;
        RECT 132.250 0.150 132.420 0.320 ;
      LAYER met1 ;
        RECT 0.000 0.000 142.700 0.480 ;
    END
  END GND
  PIN Vref
    ANTENNADIFFAREA 20.189800 ;
    PORT
      LAYER li1 ;
        RECT 61.210 43.100 79.110 43.650 ;
        RECT 78.510 41.130 79.090 43.100 ;
        RECT 78.510 41.040 79.120 41.130 ;
        RECT 78.560 37.870 79.120 41.040 ;
        RECT 78.160 35.790 79.850 37.870 ;
        RECT 120.330 34.930 121.940 37.770 ;
        RECT 120.590 31.130 121.310 34.930 ;
        RECT 120.460 30.130 121.460 31.130 ;
      LAYER mcon ;
        RECT 78.670 36.565 79.200 37.095 ;
        RECT 120.945 36.290 121.115 36.460 ;
        RECT 120.945 35.930 121.115 36.100 ;
      LAYER met1 ;
        RECT 78.160 35.790 79.850 37.870 ;
        RECT 120.330 34.930 121.940 37.770 ;
      LAYER via ;
        RECT 78.805 36.860 79.065 37.120 ;
        RECT 78.805 36.540 79.065 36.800 ;
        RECT 120.900 36.065 121.160 36.325 ;
      LAYER met2 ;
        RECT 78.160 36.670 79.850 37.870 ;
        RECT 120.330 36.670 121.940 37.770 ;
        RECT 78.160 36.020 121.940 36.670 ;
        RECT 78.160 35.790 79.850 36.020 ;
        RECT 120.330 34.930 121.940 36.020 ;
    END
  END Vref
  PIN En
    ANTENNAGATEAREA 400.000000 ;
    PORT
      LAYER li1 ;
        RECT 95.380 9.290 96.670 10.350 ;
    END
  END En
  PIN VDD
    ANTENNADIFFAREA 61.432400 ;
    PORT
      LAYER nwell ;
        RECT 83.610 61.350 113.620 66.470 ;
        RECT 83.600 60.810 113.620 61.350 ;
        RECT 83.600 59.910 113.570 60.810 ;
        RECT 83.600 39.370 113.560 59.910 ;
        RECT 83.590 37.620 113.560 39.370 ;
        RECT 93.580 37.570 113.560 37.620 ;
        RECT 103.560 37.560 113.560 37.570 ;
      LAYER li1 ;
        RECT 84.290 65.430 86.630 65.620 ;
        RECT 85.160 58.950 86.000 65.430 ;
        RECT 88.030 65.280 88.510 65.760 ;
        RECT 91.450 65.280 91.930 65.760 ;
        RECT 94.600 65.430 96.860 65.620 ;
        RECT 85.070 57.950 86.070 58.950 ;
        RECT 95.170 58.910 96.010 65.430 ;
        RECT 98.280 65.280 98.760 65.760 ;
        RECT 101.130 65.280 101.610 65.760 ;
        RECT 104.700 65.430 106.650 65.620 ;
        RECT 95.070 57.910 96.070 58.910 ;
        RECT 105.210 58.900 106.050 65.430 ;
        RECT 107.480 65.280 107.960 65.760 ;
        RECT 110.310 65.280 110.790 65.760 ;
        RECT 133.650 65.430 136.230 65.610 ;
        RECT 105.070 57.900 106.070 58.900 ;
        RECT 134.330 56.040 135.150 65.430 ;
        RECT 134.320 52.310 135.150 56.040 ;
        RECT 134.320 52.250 135.050 52.310 ;
      LAYER mcon ;
        RECT 84.305 65.435 84.475 65.605 ;
        RECT 84.965 65.435 85.135 65.605 ;
        RECT 85.745 65.435 85.915 65.605 ;
        RECT 86.445 65.435 86.615 65.605 ;
        RECT 88.185 65.430 88.355 65.600 ;
        RECT 91.605 65.430 91.775 65.600 ;
        RECT 94.605 65.435 94.775 65.605 ;
        RECT 95.345 65.435 95.515 65.605 ;
        RECT 96.105 65.435 96.275 65.605 ;
        RECT 96.685 65.435 96.855 65.605 ;
        RECT 98.435 65.430 98.605 65.600 ;
        RECT 101.285 65.430 101.455 65.600 ;
        RECT 104.715 65.435 104.885 65.605 ;
        RECT 105.315 65.435 105.485 65.605 ;
        RECT 105.945 65.435 106.115 65.605 ;
        RECT 106.475 65.435 106.645 65.605 ;
        RECT 107.635 65.430 107.805 65.600 ;
        RECT 110.465 65.430 110.635 65.600 ;
        RECT 133.665 65.435 133.835 65.605 ;
        RECT 134.515 65.435 134.685 65.605 ;
        RECT 135.245 65.435 135.415 65.605 ;
        RECT 136.055 65.435 136.225 65.605 ;
      LAYER met1 ;
        RECT 0.000 65.280 142.700 65.760 ;
    END
  END VDD
  OBS
      LAYER li1 ;
        RECT 12.840 43.610 17.640 43.710 ;
        RECT 12.840 43.160 17.660 43.610 ;
        RECT 12.840 43.080 17.640 43.160 ;
        RECT 12.880 21.650 13.380 43.080 ;
        RECT 91.120 40.010 92.120 41.010 ;
        RECT 86.200 35.230 87.320 39.130 ;
        RECT 91.270 36.110 91.990 40.010 ;
        RECT 101.080 39.910 102.080 40.910 ;
        RECT 111.030 40.850 112.030 40.900 ;
        RECT 111.030 40.820 115.280 40.850 ;
        RECT 111.030 39.990 115.310 40.820 ;
        RECT 101.200 36.700 102.010 39.910 ;
        RECT 111.030 39.900 112.030 39.990 ;
        RECT 103.100 36.750 103.910 39.180 ;
        RECT 103.100 36.700 103.940 36.750 ;
        RECT 97.900 36.310 103.940 36.700 ;
        RECT 80.440 35.220 87.320 35.230 ;
        RECT 79.600 35.210 87.320 35.220 ;
        RECT 91.260 35.550 96.640 36.110 ;
        RECT 97.840 35.770 103.940 36.310 ;
        RECT 97.840 35.740 103.800 35.770 ;
        RECT 71.930 33.780 72.650 34.460 ;
        RECT 79.600 34.350 87.300 35.210 ;
        RECT 91.260 35.200 96.660 35.550 ;
        RECT 89.410 34.390 90.480 34.730 ;
        RECT 91.270 34.390 91.940 35.200 ;
        RECT 72.130 32.160 72.500 33.780 ;
        RECT 79.600 31.310 80.440 34.350 ;
        RECT 89.410 34.250 91.940 34.390 ;
        RECT 89.410 33.690 91.910 34.250 ;
        RECT 89.410 33.380 90.480 33.690 ;
        RECT 93.520 31.990 94.480 35.200 ;
        RECT 79.530 30.310 80.530 31.310 ;
        RECT 87.310 31.220 88.310 31.280 ;
        RECT 95.850 31.270 96.660 35.200 ;
        RECT 97.840 33.940 98.800 35.740 ;
        RECT 97.850 31.270 98.760 33.940 ;
        RECT 89.740 31.220 90.740 31.270 ;
        RECT 87.310 30.350 90.740 31.220 ;
        RECT 87.310 30.280 88.310 30.350 ;
        RECT 89.740 30.270 90.740 30.350 ;
        RECT 95.740 30.270 96.740 31.270 ;
        RECT 97.790 30.270 98.790 31.270 ;
        RECT 103.800 31.160 104.800 31.230 ;
        RECT 106.240 31.160 107.240 31.270 ;
        RECT 114.500 31.170 115.310 39.990 ;
        RECT 103.800 30.320 107.240 31.160 ;
        RECT 103.800 30.230 104.800 30.320 ;
        RECT 106.240 30.270 107.240 30.320 ;
        RECT 114.410 30.170 115.410 31.170 ;
        RECT 12.660 20.960 13.500 21.650 ;
        RECT 12.625 18.055 13.415 18.845 ;
        RECT 17.495 18.055 18.285 18.845 ;
        RECT 22.715 17.945 23.505 18.735 ;
        RECT 27.585 17.945 28.375 18.735 ;
        RECT 32.685 17.945 33.475 18.735 ;
        RECT 55.200 14.980 60.460 15.010 ;
        RECT 48.070 14.960 50.280 14.970 ;
        RECT 48.050 14.400 50.280 14.960 ;
        RECT 55.180 14.400 60.460 14.980 ;
        RECT 48.070 14.390 50.280 14.400 ;
        RECT 55.200 14.370 60.460 14.400 ;
        RECT 59.180 14.050 60.430 14.370 ;
        RECT 12.505 12.925 13.295 13.715 ;
        RECT 17.725 13.075 18.515 13.865 ;
        RECT 22.745 13.015 23.535 13.805 ;
        RECT 27.595 13.015 28.385 13.805 ;
        RECT 32.685 13.075 33.475 13.865 ;
        RECT 55.760 6.410 56.280 7.110 ;
        RECT 59.180 5.360 60.460 14.050 ;
        RECT 134.330 13.990 135.070 17.710 ;
        RECT 134.350 13.770 135.010 13.990 ;
        RECT 72.540 11.970 72.870 12.300 ;
        RECT 81.300 12.270 82.300 13.270 ;
        RECT 112.270 12.310 113.270 13.310 ;
        RECT 72.570 9.190 72.850 11.970 ;
        RECT 72.260 8.280 73.030 9.190 ;
        RECT 75.790 9.010 76.460 9.320 ;
        RECT 77.470 9.010 78.500 11.340 ;
        RECT 81.490 9.720 82.040 12.270 ;
        RECT 75.790 8.520 78.500 9.010 ;
        RECT 80.720 8.560 82.140 9.720 ;
        RECT 112.550 9.450 113.030 12.310 ;
        RECT 122.960 12.300 123.960 13.300 ;
        RECT 128.950 13.190 129.950 13.290 ;
        RECT 134.370 13.190 135.010 13.770 ;
        RECT 128.950 12.380 135.030 13.190 ;
        RECT 75.790 8.270 76.460 8.520 ;
        RECT 77.470 8.060 78.500 8.520 ;
        RECT 112.290 8.460 113.280 9.450 ;
        RECT 123.090 8.130 123.820 12.300 ;
        RECT 128.950 12.290 129.950 12.380 ;
        RECT 109.770 8.060 123.820 8.130 ;
        RECT 77.470 7.330 123.820 8.060 ;
        RECT 77.470 7.320 82.020 7.330 ;
        RECT 82.460 7.320 123.820 7.330 ;
        RECT 77.470 7.270 78.500 7.320 ;
        RECT 79.200 7.280 82.020 7.320 ;
        RECT 109.290 7.270 123.820 7.320 ;
        RECT 66.470 5.360 68.780 6.030 ;
        RECT 59.120 4.000 68.780 5.360 ;
        RECT 66.470 3.450 68.780 4.000 ;
        RECT 75.010 5.360 76.440 5.880 ;
        RECT 97.830 5.380 98.770 5.410 ;
        RECT 111.760 5.380 113.530 5.580 ;
        RECT 97.380 5.370 113.530 5.380 ;
        RECT 84.590 5.360 113.530 5.370 ;
        RECT 75.010 4.220 113.530 5.360 ;
        RECT 75.010 4.210 111.950 4.220 ;
        RECT 75.010 3.640 76.440 4.210 ;
        RECT 84.590 4.200 98.980 4.210 ;
        RECT 97.380 4.180 98.980 4.200 ;
      LAYER mcon ;
        RECT 72.210 34.045 72.380 34.215 ;
        RECT 89.815 34.120 89.985 34.290 ;
        RECT 89.815 33.760 89.985 33.930 ;
        RECT 12.930 21.190 13.100 21.360 ;
        RECT 12.695 18.605 12.865 18.775 ;
        RECT 13.175 18.605 13.345 18.775 ;
        RECT 12.695 18.125 12.865 18.295 ;
        RECT 13.175 18.125 13.345 18.295 ;
        RECT 17.565 18.605 17.735 18.775 ;
        RECT 18.045 18.605 18.215 18.775 ;
        RECT 17.565 18.125 17.735 18.295 ;
        RECT 18.045 18.125 18.215 18.295 ;
        RECT 22.785 18.495 22.955 18.665 ;
        RECT 23.265 18.495 23.435 18.665 ;
        RECT 22.785 18.015 22.955 18.185 ;
        RECT 23.265 18.015 23.435 18.185 ;
        RECT 27.655 18.495 27.825 18.665 ;
        RECT 28.135 18.495 28.305 18.665 ;
        RECT 27.655 18.015 27.825 18.185 ;
        RECT 28.135 18.015 28.305 18.185 ;
        RECT 32.755 18.495 32.925 18.665 ;
        RECT 33.235 18.495 33.405 18.665 ;
        RECT 32.755 18.015 32.925 18.185 ;
        RECT 33.235 18.015 33.405 18.185 ;
        RECT 48.765 14.610 48.935 14.780 ;
        RECT 49.125 14.610 49.295 14.780 ;
        RECT 49.485 14.610 49.655 14.780 ;
        RECT 12.575 13.475 12.745 13.645 ;
        RECT 13.055 13.475 13.225 13.645 ;
        RECT 12.575 12.995 12.745 13.165 ;
        RECT 13.055 12.995 13.225 13.165 ;
        RECT 17.795 13.625 17.965 13.795 ;
        RECT 18.275 13.625 18.445 13.795 ;
        RECT 17.795 13.145 17.965 13.315 ;
        RECT 18.275 13.145 18.445 13.315 ;
        RECT 22.815 13.565 22.985 13.735 ;
        RECT 23.295 13.565 23.465 13.735 ;
        RECT 22.815 13.085 22.985 13.255 ;
        RECT 23.295 13.085 23.465 13.255 ;
        RECT 27.665 13.565 27.835 13.735 ;
        RECT 28.145 13.565 28.315 13.735 ;
        RECT 27.665 13.085 27.835 13.255 ;
        RECT 28.145 13.085 28.315 13.255 ;
        RECT 32.755 13.625 32.925 13.795 ;
        RECT 33.235 13.625 33.405 13.795 ;
        RECT 32.755 13.145 32.925 13.315 ;
        RECT 33.235 13.145 33.405 13.315 ;
        RECT 55.935 6.855 56.105 7.025 ;
        RECT 55.935 6.495 56.105 6.665 ;
        RECT 72.555 8.675 72.725 8.845 ;
        RECT 75.985 8.655 76.155 8.825 ;
        RECT 81.310 8.985 81.480 9.155 ;
        RECT 112.750 8.840 112.920 9.010 ;
        RECT 67.155 4.145 67.685 5.035 ;
        RECT 75.655 4.710 75.825 4.880 ;
        RECT 112.340 4.525 112.870 5.055 ;
        RECT 75.655 4.350 75.825 4.520 ;
      LAYER met1 ;
        RECT 71.930 33.780 72.650 34.460 ;
        RECT 89.410 33.380 90.480 34.730 ;
        RECT 12.660 20.960 13.500 21.650 ;
        RECT 12.770 18.865 13.280 20.960 ;
        RECT 12.605 18.035 13.435 18.865 ;
        RECT 17.475 18.660 18.305 18.865 ;
        RECT 22.695 18.660 23.525 18.755 ;
        RECT 27.565 18.660 28.395 18.755 ;
        RECT 32.665 18.680 33.495 18.755 ;
        RECT 32.665 18.660 49.050 18.680 ;
        RECT 17.475 18.190 49.050 18.660 ;
        RECT 17.475 18.035 18.305 18.190 ;
        RECT 17.840 13.885 18.230 18.035 ;
        RECT 22.695 17.925 23.525 18.190 ;
        RECT 27.565 17.925 28.395 18.190 ;
        RECT 32.665 18.040 49.050 18.190 ;
        RECT 32.665 17.925 33.495 18.040 ;
        RECT 46.940 18.000 49.050 18.040 ;
        RECT 48.270 15.060 49.050 18.000 ;
        RECT 48.270 14.960 50.080 15.060 ;
        RECT 48.050 14.400 50.270 14.960 ;
        RECT 12.485 13.660 13.315 13.735 ;
        RECT 17.705 13.660 18.535 13.885 ;
        RECT 22.725 13.660 23.555 13.825 ;
        RECT 27.575 13.660 28.405 13.825 ;
        RECT 12.485 13.190 28.405 13.660 ;
        RECT 12.485 12.905 13.315 13.190 ;
        RECT 17.705 13.055 18.535 13.190 ;
        RECT 22.725 12.995 23.555 13.190 ;
        RECT 27.575 12.995 28.405 13.190 ;
        RECT 32.665 13.790 33.495 13.885 ;
        RECT 32.665 13.180 45.710 13.790 ;
        RECT 32.665 13.055 33.495 13.180 ;
        RECT 45.230 6.980 45.680 13.180 ;
        RECT 72.270 9.180 72.570 9.200 ;
        RECT 72.850 9.180 73.030 9.200 ;
        RECT 72.270 8.280 73.030 9.180 ;
        RECT 75.770 9.120 76.470 9.320 ;
        RECT 75.770 8.540 76.490 9.120 ;
        RECT 80.720 8.560 82.140 9.720 ;
        RECT 112.290 9.430 112.550 9.440 ;
        RECT 113.030 9.430 113.290 9.440 ;
        RECT 75.770 8.260 76.470 8.540 ;
        RECT 112.290 8.440 113.290 9.430 ;
        RECT 55.190 6.980 56.990 8.040 ;
        RECT 45.230 6.310 56.990 6.980 ;
        RECT 45.260 6.280 56.990 6.310 ;
        RECT 55.190 5.600 56.990 6.280 ;
        RECT 66.500 5.180 68.790 6.030 ;
        RECT 66.460 4.160 68.790 5.180 ;
        RECT 66.500 3.450 68.790 4.160 ;
        RECT 75.020 5.340 76.460 5.850 ;
        RECT 111.760 5.340 113.530 5.580 ;
        RECT 75.020 4.240 76.470 5.340 ;
        RECT 111.750 4.240 113.530 5.340 ;
        RECT 75.020 3.640 76.460 4.240 ;
        RECT 111.760 4.220 113.530 4.240 ;
      LAYER via ;
        RECT 72.165 34.000 72.425 34.260 ;
        RECT 89.770 34.055 90.030 34.315 ;
        RECT 89.770 33.735 90.030 33.995 ;
        RECT 72.520 8.610 72.780 8.870 ;
        RECT 75.985 8.605 76.245 8.865 ;
        RECT 81.265 8.940 81.525 9.200 ;
        RECT 112.710 8.800 112.970 9.060 ;
        RECT 67.145 4.135 67.725 5.035 ;
        RECT 75.650 4.650 75.910 4.910 ;
        RECT 75.650 4.330 75.910 4.590 ;
        RECT 112.475 4.655 112.735 4.915 ;
      LAYER met2 ;
        RECT 71.930 34.220 72.650 34.460 ;
        RECT 89.410 34.220 90.480 34.730 ;
        RECT 71.930 33.950 90.480 34.220 ;
        RECT 71.930 33.780 72.650 33.950 ;
        RECT 79.510 33.930 80.650 33.950 ;
        RECT 89.410 33.380 90.480 33.950 ;
        RECT 72.270 9.180 72.570 9.200 ;
        RECT 72.850 9.180 73.030 9.200 ;
        RECT 72.270 9.100 73.030 9.180 ;
        RECT 75.770 9.100 76.470 9.320 ;
        RECT 72.270 8.460 76.470 9.100 ;
        RECT 80.720 8.560 82.140 9.720 ;
        RECT 112.290 9.430 112.550 9.440 ;
        RECT 113.030 9.430 113.290 9.440 ;
        RECT 72.270 8.280 73.030 8.460 ;
        RECT 73.460 8.450 74.740 8.460 ;
        RECT 75.770 8.260 76.470 8.460 ;
        RECT 55.190 7.050 56.990 8.040 ;
        RECT 81.170 7.050 81.910 8.560 ;
        RECT 112.290 8.440 113.290 9.430 ;
        RECT 55.190 6.350 81.930 7.050 ;
        RECT 112.470 6.600 112.860 8.440 ;
        RECT 55.190 5.600 56.990 6.350 ;
        RECT 81.170 6.310 81.910 6.350 ;
        RECT 66.500 5.420 68.790 6.030 ;
        RECT 71.070 5.420 71.590 5.430 ;
        RECT 75.020 5.420 76.460 5.850 ;
        RECT 112.480 5.580 112.860 6.600 ;
        RECT 66.500 3.980 76.460 5.420 ;
        RECT 111.760 4.220 113.530 5.580 ;
        RECT 66.500 3.450 68.790 3.980 ;
        RECT 75.020 3.640 76.460 3.980 ;
  END
END BGR
END LIBRARY

