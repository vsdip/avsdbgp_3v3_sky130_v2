magic
tech sky130A
timestamp 1620722909
<< mvndiff >>
rect -8 17 25 25
rect -8 0 0 17
rect 17 0 25 17
rect -8 -8 25 0
<< mvndiffc >>
rect 0 0 17 17
<< locali >>
rect -8 17 25 25
rect -8 0 0 17
rect 17 0 25 17
rect -8 -8 25 0
<< end >>
