magic
tech sky130A
magscale 1 2
timestamp 1616493613
<< nwell >>
rect 11000 2800 17600 3400
<< pwell >>
rect 9030 -8892 9166 -8464
rect -1946 -10088 2314 -8912
rect 6612 -10016 18502 -9002
<< mvndiffc >>
rect 7130 -3990 7170 -3930
rect 13240 -4060 13360 -3940
rect 13534 -4032 13660 -3920
rect 17840 -4060 17960 -3940
rect 6830 -7870 6870 -7810
rect 10530 -7862 10616 -7776
<< mvpdiffc >>
rect 11440 2240 11560 2360
rect 13640 2240 13754 2352
rect 15840 2240 15954 2352
rect 12640 -1560 12760 -1440
rect 14840 -1560 14960 -1440
rect 17040 -1560 17160 -1440
<< poly >>
rect 11600 -2000 12600 -1700
rect 13800 -2000 14800 -1700
rect 16000 -2000 17000 -1700
rect 11600 -2040 17000 -2000
rect 11600 -2160 11640 -2040
rect 11760 -2160 13640 -2040
rect 13760 -2160 15320 -2040
rect 15440 -2160 17000 -2040
rect 11600 -2200 17000 -2160
rect 7598 -3204 17802 -2800
rect 7598 -3208 13694 -3204
rect 15198 -3208 17802 -3204
rect 7600 -3802 8602 -3208
rect 10688 -3210 11802 -3208
rect 10688 -3404 11674 -3210
rect 9198 -3640 10198 -3602
rect 9198 -3780 9220 -3640
rect 9380 -3780 10198 -3640
rect 9198 -3804 10198 -3780
rect 10688 -3818 11672 -3404
rect 15198 -3802 16200 -3208
rect 16798 -3802 17800 -3208
rect 6900 -8200 7100 -8002
rect 10804 -8198 11280 -8192
rect 10356 -8200 11280 -8198
rect 12200 -8200 13202 -8000
rect 13698 -8102 14698 -7978
rect 13698 -8200 14704 -8102
rect 6898 -8240 14704 -8200
rect 6898 -8360 13240 -8240
rect 13360 -8360 14704 -8240
rect 6898 -8400 14704 -8360
rect 10356 -8402 10816 -8400
<< polycont >>
rect 11640 -2160 11760 -2040
rect 13640 -2160 13760 -2040
rect 15320 -2160 15440 -2040
rect 9220 -3780 9380 -3640
rect 13240 -8360 13360 -8240
<< locali >>
rect 11422 2360 11574 2380
rect 11422 2240 11440 2360
rect 11560 2240 11574 2360
rect 11422 2222 11574 2240
rect 13620 2352 13772 2372
rect 13620 2240 13640 2352
rect 13754 2240 13772 2352
rect 13620 2220 13772 2240
rect 15820 2352 15972 2372
rect 15820 2240 15840 2352
rect 15954 2240 15972 2352
rect 15820 2220 15972 2240
rect -134 116 362 200
rect -134 46 62 116
rect 162 46 362 116
rect -134 -38 362 46
rect 7342 112 7786 196
rect 7342 50 7478 112
rect 7622 50 7786 112
rect 7342 -16 7786 50
rect 12620 -1440 12780 -1420
rect 12620 -1560 12640 -1440
rect 12760 -1560 12780 -1440
rect 12620 -1580 12780 -1560
rect 14820 -1440 14980 -1420
rect 14820 -1560 14840 -1440
rect 14960 -1560 14980 -1440
rect 14820 -1580 14980 -1560
rect 17020 -1440 17180 -1420
rect 17020 -1560 17040 -1440
rect 17160 -1560 17180 -1440
rect 17020 -1580 17180 -1560
rect -3478 -1666 -3002 -1590
rect -3478 -1704 -3326 -1666
rect -3164 -1704 -3002 -1666
rect -3478 -1790 -3002 -1704
rect 6268 -1662 6758 -1586
rect 6268 -1736 6418 -1662
rect 6568 -1736 6758 -1662
rect 6268 -1812 6758 -1736
rect 11618 -2040 11780 -2020
rect 11618 -2160 11640 -2040
rect 11760 -2160 11780 -2040
rect 11618 -2182 11780 -2160
rect 13620 -2040 13780 -2020
rect 13620 -2160 13640 -2040
rect 13760 -2160 13780 -2040
rect 13620 -2180 13780 -2160
rect 15300 -2040 15460 -2020
rect 15300 -2160 15320 -2040
rect 15440 -2160 15460 -2040
rect 15300 -2180 15460 -2160
rect 9200 -3640 9400 -3620
rect 9200 -3780 9220 -3640
rect 9380 -3780 9400 -3640
rect 9200 -3800 9400 -3780
rect 7110 -3930 7190 -3910
rect 13508 -3920 13692 -3902
rect 7110 -3990 7130 -3930
rect 7170 -3990 7190 -3930
rect 7110 -4010 7190 -3990
rect 13220 -3940 13380 -3920
rect 13220 -4060 13240 -3940
rect 13360 -4060 13380 -3940
rect 13220 -4080 13380 -4060
rect 13508 -4032 13534 -3920
rect 13660 -4032 13692 -3920
rect 13508 -4064 13692 -4032
rect 17820 -3940 17980 -3920
rect 17820 -4060 17840 -3940
rect 17960 -4060 17980 -3940
rect 17820 -4080 17980 -4060
rect 4128 -7508 4606 -7432
rect -1020 -7582 -868 -7510
rect 4128 -7584 4302 -7508
rect 4424 -7584 4606 -7508
rect 4128 -7646 4606 -7584
rect 5650 -7516 6118 -7440
rect 5650 -7588 5810 -7516
rect 5936 -7588 6118 -7516
rect 5650 -7646 6118 -7588
rect -2452 -7864 -2024 -7812
rect -1578 -7864 -1512 -7738
rect 78 -7846 144 -7704
rect 894 -7846 960 -7704
rect 1702 -7850 1768 -7708
rect 10490 -7776 10672 -7718
rect 6806 -7810 6890 -7790
rect -2452 -7958 2092 -7864
rect 6806 -7870 6830 -7810
rect 6870 -7870 6890 -7810
rect 6806 -7890 6890 -7870
rect 10490 -7862 10530 -7776
rect 10616 -7862 10672 -7776
rect 10490 -7894 10672 -7862
rect -2452 -8024 -2300 -7958
rect -2200 -8024 2092 -7958
rect -2452 -8042 2092 -8024
rect -2452 -8116 -2024 -8042
rect 13220 -8240 13380 -8220
rect 13220 -8360 13240 -8240
rect 13360 -8360 13380 -8240
rect 13220 -8380 13380 -8360
rect -1562 -8734 -1496 -8592
rect -750 -8722 -684 -8580
rect 90 -8700 156 -8558
rect 894 -8700 960 -8558
rect 1702 -8708 1768 -8566
<< viali >>
rect 11440 2240 11560 2360
rect 13640 2240 13754 2352
rect 15840 2240 15954 2352
rect 62 46 162 116
rect 7478 50 7622 112
rect 12640 -1560 12760 -1440
rect 14840 -1560 14960 -1440
rect 17040 -1560 17160 -1440
rect -3326 -1704 -3164 -1666
rect 6418 -1736 6568 -1662
rect 11640 -2160 11760 -2040
rect 13640 -2160 13760 -2040
rect 15320 -2160 15440 -2040
rect 9220 -3780 9380 -3640
rect 7130 -3990 7170 -3930
rect 13240 -4060 13360 -3940
rect 13534 -4032 13660 -3920
rect 17840 -4060 17960 -3940
rect 4302 -7584 4424 -7508
rect 5810 -7588 5936 -7516
rect 6830 -7870 6870 -7810
rect 10530 -7862 10616 -7776
rect -2300 -8024 -2200 -7958
rect 13240 -8360 13360 -8240
<< metal1 >>
rect 11416 2360 11576 2800
rect 11416 2240 11440 2360
rect 11560 2240 11576 2360
rect 11416 2216 11576 2240
rect 13616 2352 13776 2800
rect 13616 2240 13640 2352
rect 13754 2240 13776 2352
rect 13616 2214 13776 2240
rect 15816 2352 15976 2800
rect 15816 2240 15840 2352
rect 15954 2240 15976 2352
rect 15816 2214 15976 2240
rect -134 116 362 200
rect -134 46 62 116
rect 162 46 362 116
rect -134 -38 362 46
rect 7342 112 7786 196
rect 7342 50 7478 112
rect 7622 50 7786 112
rect 7342 -16 7786 50
rect 12620 -1440 13380 -1420
rect 9502 -1580 9806 -1534
rect 12620 -1560 12640 -1440
rect 12760 -1560 13380 -1440
rect 12620 -1580 13380 -1560
rect 14820 -1440 15460 -1420
rect 14820 -1560 14840 -1440
rect 14960 -1560 15460 -1440
rect 14820 -1580 15460 -1560
rect 17020 -1440 17980 -1420
rect 17020 -1560 17040 -1440
rect 17160 -1560 17980 -1440
rect 17020 -1580 17980 -1560
rect -3478 -1666 -3002 -1590
rect -3478 -1704 -3326 -1666
rect -3164 -1704 -3002 -1666
rect -3478 -1790 -3002 -1704
rect 6268 -1636 6758 -1586
rect 7982 -1620 8474 -1610
rect 9502 -1620 9542 -1580
rect 7334 -1628 9542 -1620
rect 7158 -1636 9542 -1628
rect 6268 -1662 9542 -1636
rect 6268 -1736 6418 -1662
rect 6568 -1736 9542 -1662
rect 6268 -1778 9542 -1736
rect -3348 -7500 -3170 -1790
rect 6268 -1812 6758 -1778
rect 7158 -1780 9542 -1778
rect 7158 -1790 7366 -1780
rect 7982 -1788 8536 -1780
rect 9502 -1820 9542 -1780
rect 9760 -1820 9806 -1580
rect 9502 -1858 9806 -1820
rect 10220 -2040 11780 -2020
rect 10220 -2160 11640 -2040
rect 11760 -2160 11780 -2040
rect 10220 -2180 11780 -2160
rect 7110 -3640 9400 -3618
rect 7110 -3710 9220 -3640
rect 7110 -3930 7190 -3710
rect 8620 -3780 9220 -3710
rect 9380 -3780 9400 -3640
rect 8620 -3802 9400 -3780
rect 8620 -3924 8780 -3802
rect 10220 -3920 10380 -2180
rect 11618 -2182 11780 -2180
rect 11732 -3696 12162 -3692
rect 11732 -3798 12164 -3696
rect 7110 -3990 7130 -3930
rect 7170 -3990 7190 -3930
rect 7110 -4010 7190 -3990
rect 11734 -4012 11856 -3798
rect 12042 -4012 12164 -3798
rect 13220 -3940 13380 -1580
rect 13620 -2040 13780 -2020
rect 13620 -2160 13640 -2040
rect 13760 -2160 13780 -2040
rect 13620 -3136 13780 -2160
rect 15300 -2040 15460 -1580
rect 15300 -2160 15320 -2040
rect 15440 -2160 15460 -2040
rect 15300 -2180 15460 -2160
rect 13542 -3204 13780 -3136
rect 13542 -3478 13776 -3204
rect 13546 -3902 13678 -3478
rect 14742 -3764 15172 -3678
rect 14742 -3784 15174 -3764
rect 13220 -4060 13240 -3940
rect 13360 -4060 13380 -3940
rect 13220 -4080 13380 -4060
rect 13508 -3920 13692 -3902
rect 13508 -4032 13534 -3920
rect 13660 -4032 13692 -3920
rect 14742 -4000 14864 -3784
rect 15038 -3910 15174 -3784
rect 15038 -3924 15160 -3910
rect 17820 -3940 17980 -1580
rect 13508 -4064 13692 -4032
rect 17820 -4060 17840 -3940
rect 17960 -4060 17980 -3940
rect 17820 -4080 17980 -4060
rect 4128 -7486 4606 -7432
rect 1680 -7488 4606 -7486
rect -3348 -7586 -1576 -7500
rect -744 -7508 4606 -7488
rect -1572 -7572 -1488 -7570
rect -744 -7584 4302 -7508
rect 4424 -7584 4606 -7508
rect -3348 -7592 -1578 -7586
rect -3348 -7594 -3170 -7592
rect -744 -7598 4606 -7584
rect -2452 -7958 -2024 -7812
rect -2452 -8024 -2300 -7958
rect -2200 -8024 -2024 -7958
rect -2452 -8116 -2024 -8024
rect -3800 -9002 -2954 -9000
rect -2360 -9002 -2192 -8116
rect -742 -8350 -670 -7598
rect 1680 -7606 4606 -7598
rect 4128 -7646 4606 -7606
rect 5650 -7516 6118 -7440
rect 5650 -7588 5810 -7516
rect 5936 -7588 6118 -7516
rect 5650 -7646 6118 -7588
rect 6498 -7810 6890 -7790
rect 6498 -7870 6830 -7810
rect 6870 -7870 6890 -7810
rect 6498 -7890 6890 -7870
rect 5062 -8302 5456 -8190
rect 5062 -8344 5178 -8302
rect 4986 -8348 5178 -8344
rect -1500 -8460 934 -8350
rect 1682 -8444 5178 -8348
rect 5062 -8458 5178 -8444
rect 5332 -8458 5456 -8302
rect 5062 -8542 5456 -8458
rect 6498 -8546 6600 -7890
rect 9018 -8546 9178 -7718
rect 10490 -7776 10672 -7718
rect 10490 -7862 10530 -7776
rect 10616 -7862 10672 -7776
rect 10490 -7894 10672 -7862
rect 13222 -8220 13384 -7874
rect 13220 -8240 13384 -8220
rect 13220 -8360 13240 -8240
rect 13360 -8360 13384 -8240
rect 13220 -8380 13384 -8360
rect 6500 -8612 6600 -8546
rect 9020 -8612 9178 -8546
rect 6504 -8878 6582 -8612
rect 9030 -8878 9166 -8612
rect 6500 -9000 6600 -8878
rect 9020 -9000 9178 -8878
rect -1948 -9002 20000 -9000
rect -3800 -9998 20000 -9002
rect -3800 -10000 -2210 -9998
rect 2694 -10000 20000 -9998
<< via1 >>
rect 62 46 162 116
rect 7478 50 7622 112
rect 9542 -1820 9760 -1580
rect 7440 -4060 7560 -3940
rect 16640 -4060 16760 -3940
rect 5810 -7588 5936 -7516
rect 5178 -8458 5332 -8302
rect 10530 -7862 10616 -7776
rect 16240 -7858 16362 -7736
<< metal2 >>
rect -134 122 362 200
rect -134 34 60 122
rect 184 34 362 122
rect -134 -38 362 34
rect 7342 112 7786 196
rect 7342 50 7478 112
rect 7622 50 7786 112
rect 7342 -16 7786 50
rect 7420 -124 7578 -16
rect 7420 -3940 7580 -124
rect 9546 -1534 9762 -1524
rect 9502 -1580 9806 -1534
rect 9502 -1820 9542 -1580
rect 9760 -1820 9806 -1580
rect 9502 -1858 9806 -1820
rect 9560 -2418 9740 -1858
rect 10140 -2418 16100 -2416
rect 9560 -2580 16780 -2418
rect 9560 -2582 10610 -2580
rect 10792 -2582 15540 -2580
rect 7420 -4060 7440 -3940
rect 7560 -4060 7580 -3940
rect 7420 -4080 7580 -4060
rect 16620 -3940 16780 -2580
rect 16620 -4060 16640 -3940
rect 16760 -4060 16780 -3940
rect 16620 -4080 16780 -4060
rect 5650 -7516 6118 -7440
rect 5650 -7588 5810 -7516
rect 5936 -7588 6118 -7516
rect 5650 -7646 6118 -7588
rect 5062 -8284 5452 -8186
rect 5062 -8458 5162 -8284
rect 5336 -8458 5452 -8284
rect 5062 -8562 5452 -8458
rect 5774 -8436 6010 -7646
rect 10490 -7776 10672 -7718
rect 10490 -7862 10530 -7776
rect 10616 -7862 10672 -7776
rect 10490 -7894 10672 -7862
rect 16220 -7736 16380 -7718
rect 16220 -7858 16240 -7736
rect 16362 -7858 16380 -7736
rect 5774 -8440 6176 -8436
rect 16220 -8440 16380 -7858
rect 5774 -8444 10382 -8440
rect 10798 -8444 16380 -8440
rect 5774 -8588 16380 -8444
rect 5774 -8600 10382 -8588
rect 10798 -8600 16380 -8588
rect 5774 -8604 6176 -8600
<< via2 >>
rect 60 116 184 122
rect 60 46 62 116
rect 62 46 162 116
rect 162 46 184 116
rect 60 34 184 46
rect 5162 -8302 5336 -8284
rect 5162 -8458 5178 -8302
rect 5178 -8458 5332 -8302
rect 5332 -8458 5336 -8302
rect 10530 -7862 10616 -7776
<< metal3 >>
rect -1128 3402 -422 3404
rect -1128 3400 134 3402
rect -3800 2800 20000 3400
rect -572 2798 286 2800
rect -36 208 286 2798
rect -142 122 362 208
rect -142 34 60 122
rect 184 34 362 122
rect -142 -32 362 34
rect -134 -38 362 -32
rect 10490 -7776 10672 -7718
rect 10490 -7806 10530 -7776
rect 10488 -7862 10530 -7806
rect 10616 -7862 10672 -7776
rect 10488 -7894 10672 -7862
rect 5062 -8284 5456 -8210
rect 5062 -8458 5162 -8284
rect 5336 -8458 5456 -8284
rect 5062 -8562 5456 -8458
rect 5172 -8654 5362 -8562
rect 5182 -8698 5362 -8654
rect 10488 -8692 10650 -7894
rect 8190 -8698 10650 -8692
rect 5182 -8854 10650 -8698
rect 5182 -8860 8230 -8854
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_5
timestamp 1615375237
transform 1 0 -1922 0 1 -7956
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_0
timestamp 1615375237
transform 1 0 -1930 0 1 -8804
box 26 26 770 795
use sub2vsscontact  sub2vsscontact_9
timestamp 1615639835
transform 1 0 -1798 0 1 -10002
box 0 0 400 1000
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_6
timestamp 1615375237
transform 1 0 -1100 0 1 -7940
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_1
timestamp 1615375237
transform 1 0 -1100 0 1 -8796
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_7
timestamp 1615375237
transform 1 0 -284 0 1 -7948
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_2
timestamp 1615375237
transform 1 0 -276 0 1 -8796
box 26 26 770 795
use sub2vsscontact  sub2vsscontact_10
timestamp 1615639835
transform 1 0 -556 0 1 -10006
box 0 0 400 1000
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_9
timestamp 1615375237
transform 1 0 1334 0 1 -7934
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_8
timestamp 1615375237
transform 1 0 530 0 1 -7932
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_4
timestamp 1615375237
transform 1 0 1328 0 1 -8780
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_3
timestamp 1615375237
transform 1 0 530 0 1 -8796
box 26 26 770 795
use sub2vsscontact  sub2vsscontact_11
timestamp 1615639835
transform 1 0 658 0 1 -10002
box 0 0 400 1000
use sub2vsscontact  sub2vsscontact_12
timestamp 1615639835
transform 1 0 1894 0 1 -9986
box 0 0 400 1000
use resistor30k  resistor30k_0
timestamp 1615979809
transform 0 1 8206 -1 0 -5880
box 1560 -4060 1762 -2096
use Nmos520  Nmos520_6
timestamp 1615565174
transform 1 0 5400 0 1 -7902
box 2000 -100 3400 4100
use Nmos120  Nmos120_0
timestamp 1615566045
transform 1 0 6800 0 1 -7902
box 0 -100 400 4100
use sub2vsscontact  sub2vsscontact_0
timestamp 1615639835
transform 1 0 6802 0 1 -10002
box 0 0 400 1000
use Nmos520  Nmos520_5
timestamp 1615565174
transform 1 0 6998 0 1 -7904
box 2000 -100 3400 4100
use nmos2metal1  nmos2metal1_8
timestamp 1615594203
transform 1 0 9018 0 1 -7880
box -20 -20 180 160
use sub2vsscontact  sub2vsscontact_1
timestamp 1615639835
transform 1 0 8198 0 1 -10004
box 0 0 400 1000
use Nmos520  Nmos520_0
timestamp 1615565174
transform 1 0 8486 0 1 -7900
box 2000 -100 3400 4100
use sub2vsscontact  sub2vsscontact_2
timestamp 1615639835
transform 1 0 9600 0 1 -10002
box 0 0 400 1000
use Nmos520  Nmos520_1
timestamp 1615565174
transform 1 0 10002 0 1 -7900
box 2000 -100 3400 4100
use sub2vsscontact  sub2vsscontact_3
timestamp 1615639835
transform 1 0 11000 0 1 -10002
box 0 0 400 1000
use nmos2metal1  nmos2metal1_1
timestamp 1615594203
transform 1 0 13222 0 1 -7880
box -20 -20 180 160
use Nmos520  Nmos520_2
timestamp 1615565174
transform 1 0 11500 0 1 -7894
box 2000 -100 3400 4100
use sub2vsscontact  sub2vsscontact_4
timestamp 1615639835
transform 1 0 12400 0 1 -10004
box 0 0 400 1000
use Nmos520  Nmos520_3
timestamp 1615565174
transform 1 0 12998 0 1 -7898
box 2000 -100 3400 4100
use sub2vsscontact  sub2vsscontact_5
timestamp 1615639835
transform 1 0 13796 0 1 -10004
box 0 0 400 1000
use nmos2metal1  nmos2metal1_5
timestamp 1615594203
transform 1 0 16220 0 1 -7878
box -20 -20 180 160
use sub2vsscontact  sub2vsscontact_6
timestamp 1615639835
transform 1 0 15200 0 1 -9998
box 0 0 400 1000
use Nmos520  Nmos520_4
timestamp 1615565174
transform 1 0 14600 0 1 -7900
box 2000 -100 3400 4100
use sub2vsscontact  sub2vsscontact_7
timestamp 1615639835
transform 1 0 16598 0 1 -10000
box 0 0 400 1000
use sub2vsscontact  sub2vsscontact_8
timestamp 1615639835
transform 1 0 18000 0 1 -10000
box 0 0 400 1000
use resistor273k  resistor273k_0
timestamp 1616322141
transform 1 0 -3016 0 1 -1730
box -484 -64 9764 140
use nmos2metal1  nmos2metal1_7
timestamp 1615594203
transform 1 0 7420 0 1 -4080
box -20 -20 180 160
use nmos2metal1  nmos2metal1_3
timestamp 1615594203
transform 1 0 8620 0 1 -4080
box -20 -20 180 160
use nmos2metal1  nmos2metal1_2
timestamp 1615594203
transform 1 0 10220 0 1 -4080
box -20 -20 180 160
use Pmos520  Pmos520_0
timestamp 1615566544
transform 1 0 11400 0 1 -1600
box -400 -400 1800 4400
use nmos2metal1  nmos2metal1_10
timestamp 1615594203
transform 1 0 12020 0 1 -4080
box -20 -20 180 160
use nmos2metal1  nmos2metal1_9
timestamp 1615594203
transform 1 0 11718 0 1 -4106
box -20 -20 180 160
use Pmos520  Pmos520_1
timestamp 1615566544
transform 1 0 13600 0 1 -1600
box -400 -400 1800 4400
use nmos2metal1  nmos2metal1_12
timestamp 1615594203
transform 1 0 15018 0 1 -4068
box -20 -20 180 160
use nmos2metal1  nmos2metal1_11
timestamp 1615594203
transform 1 0 14726 0 1 -4060
box -20 -20 180 160
use Pmos520  Pmos520_2
timestamp 1615566544
transform 1 0 15800 0 1 -1600
box -400 -400 1800 4400
use nmos2metal1  nmos2metal1_4
timestamp 1615594203
transform 1 0 16620 0 1 -4080
box -20 -20 180 160
use resistor200k  resistor200k_0
timestamp 1615980034
transform 0 1 -2028 -1 0 5738
box 5548 1932 5758 9814
use vddcontact  vddcontact_0
timestamp 1615585694
transform 1 0 11300 0 1 2800
box 0 0 400 600
use vddcontact  vddcontact_1
timestamp 1615585694
transform 1 0 13500 0 1 2800
box 0 0 400 600
use pmossub2vdd  pmossub2vdd_0
timestamp 1615590023
transform 1 0 12300 0 1 2800
box 0 0 400 600
use pmossub2vdd  pmossub2vdd_1
timestamp 1615590023
transform 1 0 14500 0 1 2800
box 0 0 400 600
use vddcontact  vddcontact_2
timestamp 1615585694
transform 1 0 15700 0 1 2800
box 0 0 400 600
use pmossub2vdd  pmossub2vdd_2
timestamp 1615590023
transform 1 0 16700 0 1 2800
box 0 0 400 600
<< labels >>
rlabel poly 15626 -3234 15626 -3234 1 En
rlabel metal3 18646 3076 18646 3076 1 VDDA
rlabel metal1 18950 -9556 18950 -9556 1 VSSA
rlabel poly 12756 -2104 12756 -2104 1 C
rlabel poly 14250 -8280 14250 -8280 1 A
rlabel metal1 17898 -2664 17898 -2664 1 H
rlabel metal1 7246 -3668 7246 -3668 1 G
rlabel metal1 3012 -9578 3012 -9578 1 VSSA
flabel metal3 18638 3072 18702 3120 0 FreeSans 2400 0 0 0 VDDA
flabel metal1 19126 -9618 19126 -9618 0 FreeSans 2400 0 0 0 VSSA
flabel poly 11152 -3194 11152 -3194 0 FreeSans 1600 0 0 0 En
flabel poly 14342 -2064 14342 -2064 0 FreeSans 1600 0 0 0 C
flabel poly 12592 -8244 12592 -8244 0 FreeSans 1600 0 0 0 A
flabel metal1 17930 -1838 17930 -1838 0 FreeSans 1600 0 0 0 H
flabel metal2 7488 -628 7488 -628 0 FreeSans 1600 0 0 0 K
flabel metal1 11930 -3766 11930 -3766 0 FreeSans 1600 0 0 0 B
flabel metal1 14912 -3746 14912 -3746 0 FreeSans 1600 0 0 0 D
flabel metal3 5684 -8832 5684 -8832 0 FreeSans 1600 0 0 0 I
flabel metal1 8890 -3664 8890 -3664 0 FreeSans 1600 0 0 0 G
flabel metal1 8206 -1710 8206 -1710 0 FreeSans 1600 0 0 0 VBGP
flabel metal1 -3292 -3736 -3292 -3736 0 FreeSans 1600 0 0 0 F
flabel metal1 3144 -7572 3144 -7572 0 FreeSans 1600 0 0 0 E
flabel metal2 5872 -7952 5896 -7926 0 FreeSans 1600 0 0 0 J
<< end >>
