magic
tech sky130A
timestamp 1619696242
<< nwell >>
rect 8361 6081 11362 6647
<< mvndiffc >>
rect 7119 1214 7136 1231
rect 7262 1221 7280 1239
<< poly >>
rect 8606 3918 8781 3920
rect 8606 3905 11075 3918
rect 8606 3901 10318 3905
rect 8606 3833 8641 3901
rect 8714 3834 10318 3901
rect 10378 3834 11075 3905
rect 8714 3833 11075 3834
rect 8606 3826 11075 3833
rect 8606 3825 8783 3826
rect 9120 3825 9225 3826
rect 8606 3821 8781 3825
rect 10047 3822 10232 3826
rect 9746 3316 9914 3317
rect 9089 3315 9575 3316
rect 9685 3315 10377 3316
rect 9089 3278 10377 3315
rect 7151 3249 7252 3263
rect 7151 3227 7222 3249
rect 7239 3227 7252 3249
rect 7151 3216 7252 3227
rect 9089 3216 9370 3278
rect 9436 3216 10377 3278
rect 9089 3213 10377 3216
rect 9089 3173 9538 3213
rect 9568 3211 10377 3213
rect 9568 3209 9752 3211
rect 9906 3173 10377 3211
rect 7470 1171 7925 1195
rect 7470 1105 7923 1171
rect 7470 1053 7763 1105
rect 7830 1053 7923 1105
rect 7470 996 7923 1053
rect 7647 995 7923 996
rect 8233 1072 8721 1211
rect 8233 1070 8932 1072
rect 10738 1070 11222 1154
rect 11546 1070 12034 1204
rect 12414 1183 12882 1187
rect 12414 1070 12892 1183
rect 8233 1022 12892 1070
rect 8233 944 9565 1022
rect 9647 944 12892 1022
rect 8233 919 12892 944
rect 8233 918 12117 919
rect 12414 918 12892 919
rect 8233 913 8932 918
<< polycont >>
rect 8641 3833 8714 3901
rect 10318 3834 10378 3905
rect 7222 3227 7239 3249
rect 9370 3216 9436 3278
rect 7763 1053 7830 1105
rect 9565 944 9647 1022
<< locali >>
rect 8429 6561 8663 6562
rect 8429 6543 8430 6561
rect 8448 6543 8496 6561
rect 8514 6543 8574 6561
rect 8592 6543 8644 6561
rect 8662 6543 8663 6561
rect 9460 6561 9686 6562
rect 9478 6543 9534 6561
rect 9552 6543 9610 6561
rect 9628 6543 9668 6561
rect 10470 6561 10665 6562
rect 10470 6543 10471 6561
rect 10489 6543 10531 6561
rect 10549 6543 10594 6561
rect 10612 6543 10647 6561
rect 13365 6543 13366 6561
rect 13384 6543 13451 6561
rect 13469 6543 13524 6561
rect 13542 6543 13605 6561
rect 8516 5849 8600 6543
rect 9517 5849 9601 6543
rect 10521 5845 10605 6543
rect 13433 5604 13515 6543
rect 13432 5231 13515 5604
rect 13432 5225 13505 5231
rect 1284 4308 1764 4371
rect 6121 4310 7911 4365
rect 1288 2165 1338 4308
rect 7851 4113 7909 4310
rect 7851 4104 7912 4113
rect 7856 3787 7912 4104
rect 8620 3901 8732 3913
rect 8620 3833 8641 3901
rect 8714 3833 8732 3901
rect 7816 3712 7985 3787
rect 7816 3654 7867 3712
rect 7920 3654 7985 3712
rect 7816 3579 7985 3654
rect 8620 3523 8732 3833
rect 9127 3611 9199 4088
rect 11120 4082 11528 4085
rect 10120 3670 10201 4010
rect 11120 3999 11531 4082
rect 10310 3905 10391 3918
rect 10310 3834 10318 3905
rect 10378 3834 10391 3905
rect 10310 3675 10391 3834
rect 10310 3670 10394 3675
rect 9790 3631 10394 3670
rect 8044 3522 8732 3523
rect 7960 3521 8732 3522
rect 9126 3555 9664 3611
rect 9784 3577 10394 3631
rect 9784 3574 10380 3577
rect 7193 3429 7265 3446
rect 7193 3397 7211 3429
rect 7248 3397 7265 3429
rect 7193 3378 7265 3397
rect 7960 3435 8730 3521
rect 9126 3520 9666 3555
rect 8941 3439 9048 3473
rect 9127 3439 9194 3520
rect 7213 3249 7250 3378
rect 7213 3227 7222 3249
rect 7239 3227 7250 3249
rect 7213 3216 7250 3227
rect 7960 3050 8044 3435
rect 8941 3434 9194 3439
rect 8941 3371 8970 3434
rect 9010 3425 9194 3434
rect 9010 3371 9191 3425
rect 8941 3369 9191 3371
rect 8941 3338 9048 3369
rect 9352 3278 9448 3520
rect 9352 3216 9370 3278
rect 9436 3216 9448 3278
rect 9352 3199 9448 3216
rect 8766 3035 9007 3122
rect 9585 3085 9666 3520
rect 9784 3394 9880 3574
rect 9785 3086 9876 3394
rect 10418 3032 10687 3116
rect 11450 3031 11531 3999
rect 12033 3647 12194 3777
rect 12033 3592 12082 3647
rect 12124 3592 12194 3647
rect 12033 3493 12194 3592
rect 12059 3077 12131 3493
rect 1266 2137 1350 2165
rect 1266 2118 1289 2137
rect 1314 2118 1350 2137
rect 1266 2096 1350 2118
rect 1275 1689 1325 1756
rect 1762 1689 1812 1756
rect 2291 1675 2341 1742
rect 2772 1679 2822 1746
rect 3289 1681 3337 1743
rect 2895 1664 3486 1667
rect 1107 1652 3486 1664
rect 541 1649 3486 1652
rect 434 1645 3486 1649
rect 405 1502 3486 1645
rect 405 1492 592 1502
rect 1107 1500 3486 1502
rect 405 284 557 1492
rect 1268 1426 1318 1493
rect 1787 1434 1837 1500
rect 2295 1426 2345 1493
rect 2783 1432 2833 1499
rect 2895 1484 3486 1500
rect 3289 1435 3337 1484
rect 4805 1482 5027 1496
rect 4805 1457 4872 1482
rect 4970 1457 5027 1482
rect 4805 1440 5027 1457
rect 5520 1437 6046 1501
rect 5918 1405 6043 1437
rect 5918 536 6046 1405
rect 13433 1399 13507 1771
rect 13435 1377 13501 1399
rect 13437 1319 13501 1377
rect 7257 1239 7284 1247
rect 7113 1231 7142 1239
rect 7113 1214 7119 1231
rect 7136 1214 7142 1231
rect 7113 1179 7142 1214
rect 7111 1175 7142 1179
rect 7257 1221 7262 1239
rect 7280 1221 7284 1239
rect 7257 1191 7284 1221
rect 6647 536 6878 603
rect 7111 594 7140 1175
rect 7257 919 7285 1191
rect 7226 899 7303 919
rect 7226 853 7242 899
rect 7286 853 7303 899
rect 7226 828 7303 853
rect 5912 520 6878 536
rect 5912 400 6700 520
rect 6647 398 6700 400
rect 6784 398 6878 520
rect 6647 345 6878 398
rect 7112 359 7140 594
rect 7354 746 7442 1288
rect 7747 1105 7850 1134
rect 7747 1053 7763 1105
rect 7830 1053 7850 1105
rect 7579 901 7646 932
rect 7747 901 7850 1053
rect 8149 972 8204 1264
rect 9538 1022 9667 1035
rect 7579 894 7850 901
rect 7579 854 7592 894
rect 7622 854 7850 894
rect 8072 923 8214 972
rect 9538 944 9565 1022
rect 9647 944 9667 1022
rect 11255 945 11303 1270
rect 9538 929 9667 944
rect 8072 891 8120 923
rect 8159 891 8214 923
rect 8072 856 8214 891
rect 11229 908 11328 945
rect 11229 877 11266 908
rect 11301 877 11328 908
rect 7579 852 7850 854
rect 7579 827 7646 852
rect 7747 806 7850 852
rect 11229 846 11328 877
rect 12309 813 12382 1318
rect 12927 1238 13503 1319
rect 10977 806 12382 813
rect 7112 335 7143 359
rect 402 33 558 284
rect 7115 33 7143 335
rect 7354 306 7444 746
rect 7747 733 12382 806
rect 7747 732 8202 733
rect 8246 732 12382 733
rect 7747 727 7850 732
rect 7920 728 8202 732
rect 10929 727 12382 732
rect 7501 536 7644 588
rect 9783 538 9877 541
rect 11176 538 11353 558
rect 9738 537 11353 538
rect 8459 536 11353 537
rect 7501 506 11353 536
rect 7501 500 11234 506
rect 7501 423 7548 500
rect 7600 452 11234 500
rect 11287 452 11353 506
rect 7600 423 11353 452
rect 7501 422 11353 423
rect 7501 421 11195 422
rect 7501 364 7644 421
rect 8459 420 9898 421
rect 9738 418 9898 420
rect 7355 33 7441 306
rect 353 15 380 33
rect 398 15 425 33
rect 443 15 470 33
rect 488 15 515 33
rect 533 15 560 33
rect 578 15 605 33
rect 7008 15 7070 33
rect 7088 15 7115 33
rect 7133 15 7160 33
rect 7178 15 7266 33
rect 7283 15 7341 33
rect 7358 15 7385 33
rect 7403 15 7430 33
rect 7447 15 7535 33
rect 7583 15 7836 33
rect 7857 15 8110 33
rect 8158 15 13211 33
<< viali >>
rect 8430 6543 8448 6561
rect 8496 6543 8514 6561
rect 8574 6543 8592 6561
rect 8644 6543 8662 6561
rect 9460 6543 9478 6561
rect 9534 6543 9552 6561
rect 9610 6543 9628 6561
rect 9668 6543 9686 6561
rect 10471 6543 10489 6561
rect 10531 6543 10549 6561
rect 10594 6543 10612 6561
rect 10647 6543 10665 6561
rect 13366 6543 13384 6561
rect 13451 6543 13469 6561
rect 13524 6543 13542 6561
rect 13605 6543 13623 6561
rect 7867 3654 7920 3712
rect 7211 3397 7248 3429
rect 8970 3371 9010 3434
rect 12082 3592 12124 3647
rect 1289 2118 1314 2137
rect 4872 1457 4970 1482
rect 5576 641 5628 711
rect 7242 853 7286 899
rect 6700 398 6784 520
rect 7592 854 7622 894
rect 8120 891 8159 923
rect 11266 877 11301 908
rect 7548 423 7600 500
rect 11234 452 11287 506
rect 335 15 353 33
rect 380 15 398 33
rect 425 15 443 33
rect 470 15 488 33
rect 515 15 533 33
rect 560 15 578 33
rect 605 15 623 33
rect 7070 15 7088 33
rect 7115 15 7133 33
rect 7160 15 7178 33
rect 7341 15 7358 33
rect 7385 15 7403 33
rect 7430 15 7447 33
<< metal1 >>
rect 0 6561 14270 6576
rect 0 6543 8430 6561
rect 8448 6543 8496 6561
rect 8514 6543 8574 6561
rect 8592 6543 8644 6561
rect 8662 6543 9460 6561
rect 9478 6543 9534 6561
rect 9552 6543 9610 6561
rect 9628 6543 9668 6561
rect 9686 6543 10471 6561
rect 10489 6543 10531 6561
rect 10549 6543 10594 6561
rect 10612 6543 10647 6561
rect 10665 6543 13366 6561
rect 13384 6543 13451 6561
rect 13469 6543 13524 6561
rect 13542 6543 13605 6561
rect 13623 6543 14270 6561
rect 0 6528 14270 6543
rect 7816 3712 7985 3787
rect 7816 3654 7867 3712
rect 7920 3654 7985 3712
rect 7816 3579 7985 3654
rect 12033 3647 12194 3777
rect 12033 3592 12082 3647
rect 12124 3592 12194 3647
rect 12033 3493 12194 3592
rect 7193 3429 7265 3446
rect 7193 3397 7211 3429
rect 7248 3397 7265 3429
rect 7193 3378 7265 3397
rect 8941 3434 9048 3473
rect 8941 3371 8970 3434
rect 9010 3371 9048 3434
rect 8941 3338 9048 3371
rect 1266 2137 1350 2165
rect 1266 2118 1289 2137
rect 1314 2118 1350 2137
rect 1266 2096 1350 2118
rect 1277 1834 1328 2096
rect 3282 1866 4905 1868
rect 1758 1819 4905 1866
rect 1784 1366 1823 1819
rect 3282 1804 4905 1819
rect 4694 1800 4905 1804
rect 4827 1506 4905 1800
rect 4827 1496 5008 1506
rect 4805 1482 5027 1496
rect 4805 1457 4872 1482
rect 4970 1457 5027 1482
rect 4805 1440 5027 1457
rect 1259 1319 2784 1366
rect 3277 1318 4571 1379
rect 4523 698 4568 1318
rect 7227 918 7257 920
rect 7285 918 7303 920
rect 7227 899 7303 918
rect 7227 853 7242 899
rect 7286 853 7303 899
rect 7227 852 7245 853
rect 7285 852 7303 853
rect 7227 828 7303 852
rect 7577 912 7647 932
rect 8072 923 8214 972
rect 7577 894 7649 912
rect 7577 854 7592 894
rect 7622 893 7649 894
rect 7626 854 7649 893
rect 8072 891 8120 923
rect 8159 891 8214 923
rect 8072 856 8214 891
rect 11229 943 11255 944
rect 11303 943 11329 944
rect 11229 908 11329 943
rect 11229 878 11265 908
rect 11303 878 11329 908
rect 11229 877 11266 878
rect 11301 877 11329 878
rect 7577 826 7647 854
rect 11229 844 11329 877
rect 5519 711 5699 804
rect 5519 698 5576 711
rect 4523 641 5576 698
rect 5628 641 5699 711
rect 4523 631 5699 641
rect 4526 628 5699 631
rect 5519 560 5699 628
rect 6650 520 6879 603
rect 6650 518 6700 520
rect 6784 518 6879 520
rect 6646 416 6700 518
rect 6650 398 6700 416
rect 6786 399 6879 518
rect 6784 398 6879 399
rect 6650 345 6879 398
rect 7502 534 7646 585
rect 11176 534 11353 558
rect 7502 500 7647 534
rect 7502 423 7548 500
rect 7603 424 7647 500
rect 11175 507 11353 534
rect 11175 450 11234 507
rect 11287 450 11353 507
rect 11175 424 11353 450
rect 7600 423 7646 424
rect 7502 364 7646 423
rect 11176 422 11353 424
rect 0 33 14270 48
rect 0 15 335 33
rect 353 15 380 33
rect 398 15 425 33
rect 443 15 470 33
rect 488 15 515 33
rect 533 15 560 33
rect 578 15 605 33
rect 623 15 7070 33
rect 7088 15 7115 33
rect 7133 15 7160 33
rect 7178 15 7341 33
rect 7358 15 7385 33
rect 7403 15 7430 33
rect 7447 15 14270 33
rect 0 0 14270 15
<< via1 >>
rect 7867 3654 7920 3712
rect 12082 3592 12124 3647
rect 7211 3397 7248 3429
rect 8970 3371 9010 3434
rect 7245 853 7285 896
rect 7245 852 7285 853
rect 7597 854 7622 893
rect 7622 854 7626 893
rect 8120 891 8159 923
rect 11265 878 11266 908
rect 11266 878 11301 908
rect 11301 878 11303 908
rect 6701 399 6784 518
rect 6784 399 6786 518
rect 7553 424 7600 500
rect 7600 424 7603 500
rect 11234 506 11287 507
rect 11234 452 11287 506
rect 11234 450 11287 452
<< metal2 >>
rect 7816 3712 7985 3787
rect 7816 3654 7867 3712
rect 7920 3667 7985 3712
rect 12033 3667 12194 3777
rect 7920 3654 12194 3667
rect 7816 3647 12194 3654
rect 7816 3602 12082 3647
rect 7816 3579 7985 3602
rect 12033 3592 12082 3602
rect 12124 3592 12194 3647
rect 12033 3493 12194 3592
rect 7193 3429 7265 3446
rect 7193 3397 7211 3429
rect 7248 3422 7265 3429
rect 8941 3434 9048 3473
rect 8941 3422 8970 3434
rect 7248 3397 8970 3422
rect 7193 3395 8970 3397
rect 7193 3378 7265 3395
rect 7951 3393 8065 3395
rect 8941 3371 8970 3395
rect 9010 3371 9048 3434
rect 8941 3338 9048 3371
rect 7227 918 7257 920
rect 7285 918 7303 920
rect 7227 910 7303 918
rect 7577 910 7647 932
rect 7227 896 7647 910
rect 7227 852 7245 896
rect 7285 893 7647 896
rect 7285 854 7597 893
rect 7626 854 7647 893
rect 8072 923 8214 972
rect 8072 891 8120 923
rect 8159 891 8214 923
rect 8072 856 8214 891
rect 11229 943 11255 944
rect 11303 943 11329 944
rect 11229 908 11329 943
rect 11229 878 11265 908
rect 11303 878 11329 908
rect 7285 852 7647 854
rect 7227 846 7647 852
rect 7227 828 7303 846
rect 7346 845 7474 846
rect 7577 826 7647 846
rect 5519 705 5699 804
rect 8117 705 8191 856
rect 11229 844 11329 878
rect 5519 635 8193 705
rect 11247 660 11286 844
rect 5519 560 5699 635
rect 8117 631 8191 635
rect 6650 542 6879 603
rect 7107 542 7159 543
rect 7502 542 7646 585
rect 11248 558 11286 660
rect 6650 518 7646 542
rect 6650 399 6701 518
rect 6786 500 7646 518
rect 6786 424 7553 500
rect 7603 424 7646 500
rect 6786 399 7646 424
rect 11176 507 11353 558
rect 11176 450 11234 507
rect 11287 450 11353 507
rect 11176 422 11353 450
rect 6650 398 7646 399
rect 6650 345 6879 398
rect 7502 364 7646 398
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_0
timestamp 1619696242
transform 1 0 1091 0 1 1133
box 0 0 398 398
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_1
timestamp 1619696242
transform 1 0 1613 0 1 1148
box 0 0 398 398
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_5
timestamp 1619696242
transform 1 0 1103 0 1 1646
box 0 0 398 398
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_6
timestamp 1619696242
transform 1 0 1590 0 1 1646
box 0 0 398 398
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_2
timestamp 1619696242
transform 1 0 2115 0 1 1142
box 0 0 398 398
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_3
timestamp 1619696242
transform 1 0 2600 0 1 1142
box 0 0 398 398
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_7
timestamp 1619696242
transform 1 0 2112 0 1 1635
box 0 0 398 398
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_8
timestamp 1619696242
transform 1 0 2599 0 1 1635
box 0 0 398 398
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_4
timestamp 1619696242
transform 1 0 3109 0 1 1148
box 0 0 398 398
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_9
timestamp 1619696242
transform 1 0 3109 0 1 1635
box 0 0 398 398
use resistor30K  resistor30K_0
timestamp 1618573301
transform 1 0 5008 0 1 1450
box -201 -11 731 48
use resistor273K  resistor273K_0
timestamp 1619682155
transform 1 0 1761 0 1 4321
box -215 -5 4585 40
use nmos_substrate  nmos_substrate_3
timestamp 1619685304
transform 1 0 7810 0 1 0
box 0 0 48 48
use nmos_substrate  nmos_substrate_2
timestamp 1619685304
transform 1 0 7535 0 1 0
box 0 0 48 48
use nmos_substrate  nmos_substrate_1
timestamp 1619685304
transform 1 0 6960 0 1 0
box 0 0 48 48
use nmos_substrate  nmos_substrate_0
timestamp 1619685304
transform 1 0 7235 0 1 0
box 0 0 48 48
use NMOS520  NMOS520_0
timestamp 1618661393
transform 1 0 7455 0 1 1180
box -101 -50 601 2050
use NMOS120  NMOS120_0
timestamp 1618661559
transform 1 0 7151 0 1 1190
box -40 -30 140 2030
use nmos2metal  nmos2metal_9
timestamp 1619503262
transform 1 0 7354 0 1 1228
box 0 0 100 100
use nmos_substrate  nmos_substrate_6
timestamp 1619685304
transform 1 0 8710 0 1 0
box 0 0 48 48
use nmos_substrate  nmos_substrate_5
timestamp 1619685304
transform 1 0 8410 0 1 0
box 0 0 48 48
use nmos_substrate  nmos_substrate_4
timestamp 1619685304
transform 1 0 8110 0 1 0
box 0 0 48 48
use NMOS520  NMOS520_1
timestamp 1618661393
transform 1 0 8229 0 1 1175
box -101 -50 601 2050
use nmos2metal  nmos2metal_14
timestamp 1619503262
transform 1 0 8130 0 1 1227
box 0 0 100 100
use nmos_substrate  nmos_substrate_7
timestamp 1619685304
transform 1 0 9010 0 1 0
box 0 0 48 48
use NMOS520  NMOS520_2
timestamp 1618661393
transform 1 0 9075 0 1 1175
box -101 -50 601 2050
use NMOS520  NMOS520_3
timestamp 1618661393
transform 1 0 9879 0 1 1175
box -101 -50 601 2050
use nmos_substrate  nmos_substrate_8
timestamp 1619685304
transform 1 0 9310 0 1 0
box 0 0 48 48
use nmos_substrate  nmos_substrate_9
timestamp 1619685304
transform 1 0 9610 0 1 0
box 0 0 48 48
use NMOS520  NMOS520_4
timestamp 1618661393
transform 1 0 10723 0 1 1180
box -101 -50 601 2050
use nmos_substrate  nmos_substrate_10
timestamp 1619685304
transform 1 0 9910 0 1 0
box 0 0 48 48
use nmos_substrate  nmos_substrate_11
timestamp 1619685304
transform 1 0 10210 0 1 0
box 0 0 48 48
use nmos_substrate  nmos_substrate_12
timestamp 1619685304
transform 1 0 10510 0 1 0
box 0 0 48 48
use PMOS520  PMOS520_0
timestamp 1619510475
transform 1 0 8610 0 1 3948
box -251 -186 750 2187
use nmos2metal  nmos2metal_8
timestamp 1619503262
transform 1 0 7953 0 1 3031
box 0 0 100 100
use nmos2metal  nmos2metal_3
timestamp 1619503262
transform 1 0 8731 0 1 3028
box 0 0 100 100
use pmos2metal  pmos2metal_3
timestamp 1619503365
transform 1 0 9112 0 1 4001
box -23 -23 123 123
use nmos2metal  nmos2metal_2
timestamp 1619503262
transform 1 0 8974 0 1 3027
box 0 0 100 100
use nmos2metal  nmos2metal_1
timestamp 1619503262
transform 1 0 9779 0 1 3027
box 0 0 100 100
use nmos2metal  nmos2metal_0
timestamp 1619503262
transform 1 0 9574 0 1 3027
box 0 0 100 100
use PMOS520  PMOS520_1
timestamp 1619510475
transform 1 0 9609 0 1 3943
box -251 -186 750 2187
use pmos2metal  pmos2metal_4
timestamp 1619503365
transform 1 0 10108 0 1 3991
box -23 -23 123 123
use nmos2metal  nmos2metal_5
timestamp 1619503262
transform 1 0 10624 0 1 3027
box 0 0 100 100
use nmos2metal  nmos2metal_4
timestamp 1619503262
transform 1 0 10380 0 1 3023
box 0 0 100 100
use PMOS520  PMOS520_2
timestamp 1619510475
transform 1 0 10607 0 1 3942
box -251 -186 750 2187
use pmos_substrate  pmos_substrate_0
timestamp 1619685549
transform 1 0 8803 0 1 6528
box -33 -34 81 81
use pmos2metal  pmos2metal_0
timestamp 1619503365
transform 1 0 8507 0 1 5795
box -23 -23 123 123
use pmos_substrate  pmos_substrate_1
timestamp 1619685549
transform 1 0 9145 0 1 6528
box -33 -34 81 81
use pmos_substrate  pmos_substrate_2
timestamp 1619685549
transform 1 0 9828 0 1 6528
box -33 -34 81 81
use pmos2metal  pmos2metal_1
timestamp 1619503365
transform 1 0 9507 0 1 5791
box -23 -23 123 123
use pmos_substrate  pmos_substrate_3
timestamp 1619685549
transform 1 0 10113 0 1 6528
box -33 -34 81 81
use pmos2metal  pmos2metal_2
timestamp 1619503365
transform 1 0 10507 0 1 5790
box -23 -23 123 123
use pmos_substrate  pmos_substrate_4
timestamp 1619685549
transform 1 0 10748 0 1 6528
box -33 -34 81 81
use pmos_substrate  pmos_substrate_5
timestamp 1619685549
transform 1 0 11031 0 1 6528
box -33 -34 81 81
use nmos_substrate  nmos_substrate_13
timestamp 1619685304
transform 1 0 10810 0 1 0
box 0 0 48 48
use nmos_substrate  nmos_substrate_14
timestamp 1619685304
transform 1 0 11109 0 1 0
box 0 0 48 48
use nmos2metal  nmos2metal_11
timestamp 1619503262
transform 1 0 11227 0 1 1231
box 0 0 100 100
use pmos2metal  pmos2metal_5
timestamp 1619503365
transform 1 0 11103 0 1 3990
box -23 -23 123 123
use nmos_substrate  nmos_substrate_17
timestamp 1619685304
transform 1 0 12010 0 1 0
box 0 0 48 48
use nmos_substrate  nmos_substrate_16
timestamp 1619685304
transform 1 0 11710 0 1 0
box 0 0 48 48
use nmos_substrate  nmos_substrate_15
timestamp 1619685304
transform 1 0 11410 0 1 0
box 0 0 48 48
use NMOS520  NMOS520_5
timestamp 1618661393
transform 1 0 11544 0 1 1175
box -101 -50 601 2050
use nmos2metal  nmos2metal_6
timestamp 1619503262
transform 1 0 11441 0 1 3017
box 0 0 100 100
use nmos2metal  nmos2metal_13
timestamp 1619503262
transform 1 0 12046 0 1 3013
box 0 0 100 100
use nmos_substrate  nmos_substrate_18
timestamp 1619685304
transform 1 0 12310 0 1 0
box 0 0 48 48
use NMOS520  NMOS520_6
timestamp 1618661393
transform 1 0 12394 0 1 1180
box -101 -50 601 2050
use nmos_substrate  nmos_substrate_19
timestamp 1619685304
transform 1 0 12610 0 1 0
box 0 0 48 48
use nmos2metal  nmos2metal_10
timestamp 1619503262
transform 1 0 12296 0 1 1230
box 0 0 100 100
use nmos_substrate  nmos_substrate_21
timestamp 1619685304
transform 1 0 13210 0 1 0
box 0 0 48 48
use nmos_substrate  nmos_substrate_20
timestamp 1619685304
transform 1 0 12910 0 1 0
box 0 0 48 48
use nmos2metal  nmos2metal_7
timestamp 1619503262
transform 1 0 12895 0 1 1229
box 0 0 100 100
use resistor200K  resistor200K_0
timestamp 1618573519
transform 0 1 13455 -1 0 5253
box -350 -20 3852 51
<< labels >>
flabel space 7131 1400 7179 1579 0 FreeSans 800 0 0 0 XM10
flabel poly 9968 3185 10079 3312 0 FreeSans 800 0 0 0 A
flabel space 10507 3079 10618 3206 0 FreeSans 400 0 0 0 D
flabel space 8865 3058 8976 3185 0 FreeSans 400 0 0 0 B
flabel space 9463 3839 9574 3966 0 FreeSans 800 0 0 0 C
flabel space 11688 2209 11736 2388 0 FreeSans 1600 0 0 0 XM13
flabel space 12605 2209 12653 2388 0 FreeSans 1600 0 0 0 XM14
flabel space 7583 2162 7817 2443 0 FreeSans 1600 0 0 0 XM9
flabel space 10832 2317 11066 2598 0 FreeSans 1600 0 0 0 XM12
flabel space 8297 2150 8531 2431 0 FreeSans 1600 0 0 0 XM11
flabel space 9975 2269 10209 2550 0 FreeSans 1600 0 0 0 XM5
flabel space 9202 2281 9436 2562 0 FreeSans 1600 0 0 0 XM4
flabel space 10740 4805 10974 5086 0 FreeSans 1600 0 0 0 XM3
flabel space 9718 4757 9952 5038 0 FreeSans 1600 0 0 0 XM2
flabel space 8744 4710 8978 4991 0 FreeSans 1600 0 0 0 XM1
flabel metal1 4038 1852 4038 1852 0 FreeSans 800 0 0 0 E
rlabel poly 10618 3863 10618 3863 1 C
flabel locali 11485 3811 11485 3811 0 FreeSans 800 0 0 0 H
rlabel poly 10138 3228 10138 3228 1 A
rlabel poly 9326 3854 9326 3854 1 C
rlabel locali 8909 3066 8909 3066 1 B
rlabel locali 10565 3066 10565 3066 1 D
rlabel locali 5957 1238 5957 1238 1 J
rlabel metal1 4357 1829 4357 1829 1 E
rlabel metal1 4186 1343 4186 1343 1 I
rlabel locali 13255 1263 13255 1263 1 K
rlabel locali 10766 762 10766 762 1 G
rlabel locali 1315 2819 1315 2819 1 F
flabel metal1 5601 18 5601 18 0 FreeSans 800 0 0 0 GND
port 1 nsew
flabel locali 6646 4335 6646 4335 0 FreeSans 800 0 0 0 Vref
port 2 nsew
flabel polycont 9565 944 9647 1022 0 FreeSans 800 0 0 0 En
port 3 nsew
<< properties >>
string LEFclass CORE
string FIXED_BBOX 0 24 14270 6552
<< end >>
