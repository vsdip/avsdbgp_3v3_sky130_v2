magic
tech sky130A
timestamp 1619685549
<< nwell >>
rect -33 -34 81 81
<< mvnsubdiff >>
rect 0 35 48 48
rect 0 12 13 35
rect 35 12 48 35
rect 0 0 48 12
<< mvnsubdiffcont >>
rect 13 12 35 35
<< locali >>
rect 0 35 48 48
rect 0 12 13 35
rect 35 12 48 35
rect 0 0 48 12
<< viali >>
rect 13 12 35 35
<< metal1 >>
rect 0 35 48 48
rect 0 12 13 35
rect 35 12 48 35
rect 0 0 48 12
<< end >>
